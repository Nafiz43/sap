CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
28 D:\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
297
13 Logic Switch~
5 1729 401 0 10 11
0 96 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9365 0 0
2
43749 0
0
13 Logic Switch~
5 1900 498 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3251 0 0
2
43749 1
0
13 Logic Switch~
5 1926 457 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 V1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5481 0 0
2
43749 2
0
13 Logic Switch~
5 1817 1001 0 1 11
0 65
0
0 0 20832 180
2 0V
-7 -16 7 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7788 0 0
2
43749 3
0
13 Logic Switch~
5 1837 942 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 20832 180
2 5V
-7 -16 7 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3273 0 0
2
43749 4
0
13 Logic Switch~
5 1837 866 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 20832 180
2 5V
-7 -16 7 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3761 0 0
2
43749 5
0
13 Logic Switch~
5 1837 900 0 1 11
0 67
0
0 0 20832 180
2 0V
-7 -16 7 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3226 0 0
2
43749 6
0
13 Logic Switch~
5 142 768 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 20832 90
2 5V
11 -5 25 3
3 V27
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4244 0 0
2
5.89911e-315 5.26354e-315
0
13 Logic Switch~
5 626 571 0 1 11
0 82
0
0 0 20832 782
2 0V
-6 -21 8 -13
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5225 0 0
2
5.89911e-315 5.30499e-315
0
13 Logic Switch~
5 248 262 0 1 11
0 102
0
0 0 20832 0
2 0V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
768 0 0
2
43749 7
0
13 Logic Switch~
5 1057 1528 0 10 11
0 97 0 0 0 0 0 0 0 0
1
0
0 0 20832 0
2 5V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5735 0 0
2
43749 8
0
13 Logic Switch~
5 89 67 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 20832 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5881 0 0
2
43749 9
0
14 Logic Display~
6 1625 166 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L43
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3275 0 0
2
5.89911e-315 0
0
14 Logic Display~
6 1598 169 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L39
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4203 0 0
2
5.89911e-315 0
0
14 Logic Display~
6 1567 168 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L34
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.89911e-315 0
0
14 Logic Display~
6 1531 166 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L33
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9102 0 0
2
5.89911e-315 0
0
8 2-In OR~
219 2271 2603 0 3 22
0 21 5 20
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U23D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
5586 0 0
2
5.89911e-315 5.32571e-315
0
7 Ground~
168 1883 422 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
525 0 0
2
5.89911e-315 5.34643e-315
0
7 Ground~
168 1789 498 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6206 0 0
2
5.89911e-315 5.3568e-315
0
14 Logic Display~
6 1485 657 0 1 2
10 28
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L21
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3418 0 0
2
5.89911e-315 5.36716e-315
0
14 Logic Display~
6 1483 686 0 1 2
10 29
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L15
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9312 0 0
2
5.89911e-315 5.37752e-315
0
14 Logic Display~
6 1451 636 0 1 2
10 31
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L44
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7419 0 0
2
5.89911e-315 5.38788e-315
0
14 Logic Display~
6 1450 599 0 1 2
10 32
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L42
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
472 0 0
2
5.89911e-315 5.39306e-315
0
14 Logic Display~
6 1530 501 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L41
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4714 0 0
2
5.89911e-315 5.39824e-315
0
9 Inverter~
13 2336 2200 0 2 22
0 36 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U27A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
9386 0 0
2
5.89911e-315 5.40342e-315
0
9 Inverter~
13 2518 2693 0 2 22
0 37 9
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U26F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
7610 0 0
2
5.89911e-315 5.4086e-315
0
14 Logic Display~
6 1055 1945 0 1 2
10 41
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
43749 10
0
14 Logic Display~
6 1053 1901 0 1 2
10 43
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L20
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3608 0 0
2
43749 11
0
14 Logic Display~
6 1052 1858 0 1 2
10 38
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L19
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6397 0 0
2
43749 12
0
14 Logic Display~
6 1052 1833 0 1 2
10 42
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L18
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3967 0 0
2
43749 13
0
14 Logic Display~
6 1050 1802 0 1 2
10 44
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L17
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8621 0 0
2
43749 14
0
14 Logic Display~
6 1040 1772 0 1 2
10 45
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L16
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
43749 15
0
9 Inverter~
13 991 1949 0 2 22
0 46 41
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U26E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
7385 0 0
2
43749 16
0
9 Inverter~
13 992 1905 0 2 22
0 47 43
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U26D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
6519 0 0
2
43749 17
0
9 Inverter~
13 1002 1861 0 2 22
0 48 38
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U26C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
552 0 0
2
43749 18
0
9 Inverter~
13 1001 1836 0 2 22
0 49 42
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U26B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
5551 0 0
2
43749 19
0
9 Inverter~
13 962 1805 0 2 22
0 50 44
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U26A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
8715 0 0
2
43749 20
0
9 Inverter~
13 958 1775 0 2 22
0 51 45
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U21F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
9763 0 0
2
43749 21
0
14 Logic Display~
6 2489 2718 0 1 2
10 37
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8443 0 0
2
43749 22
0
14 Logic Display~
6 2398 2691 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L38
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3719 0 0
2
43749 23
0
14 Logic Display~
6 2372 2686 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L37
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8671 0 0
2
43749 24
0
14 Logic Display~
6 2431 2691 0 1 2
10 37
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L36
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
43749 25
0
14 Logic Display~
6 2338 2688 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L35
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
49 0 0
2
43749 26
0
14 Logic Display~
6 2158 2695 0 1 2
10 36
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L32
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6536 0 0
2
43749 27
0
14 Logic Display~
6 2072 2700 0 1 2
10 4
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L31
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3931 0 0
2
43749 28
0
14 Logic Display~
6 1968 2698 0 1 2
10 33
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L30
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4390 0 0
2
43749 29
0
14 Logic Display~
6 1838 2696 0 1 2
10 12
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L29
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3242 0 0
2
43749 30
0
14 Logic Display~
6 1690 2692 0 1 2
10 3
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L28
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6760 0 0
2
43749 31
0
14 Logic Display~
6 1494 2706 0 1 2
10 11
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L27
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5760 0 0
2
43749 32
0
14 Logic Display~
6 1358 2722 0 1 2
10 13
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L26
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3781 0 0
2
43749 33
0
14 Logic Display~
6 1259 2576 0 1 2
10 8
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L25
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8545 0 0
2
43749 34
0
14 Logic Display~
6 1163 2508 0 1 2
10 10
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L24
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9739 0 0
2
43749 35
0
14 Logic Display~
6 1099 2747 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L23
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
388 0 0
2
43749 36
0
8 2-In OR~
219 2140 2543 0 3 22
0 36 52 4
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U23B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4595 0 0
2
43749 37
0
9 2-In AND~
219 2094 2160 0 3 22
0 41 40 36
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U25B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3173 0 0
2
43749 38
0
9 Inverter~
13 2061 2553 0 2 22
0 52 33
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U21E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
9261 0 0
2
43749 39
0
9 Inverter~
13 1921 2546 0 2 22
0 53 12
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U21D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
3494 0 0
2
43749 40
0
9 2-In AND~
219 2065 2478 0 3 22
0 40 42 52
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U25A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9101 0 0
2
43749 41
0
8 2-In OR~
219 1923 2497 0 3 22
0 54 37 53
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U23A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
358 0 0
2
43749 42
0
9 2-In AND~
219 1910 2393 0 3 22
0 43 40 37
0
0 0 608 270
5 74F08
-18 -24 17 -16
4 U19B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3726 0 0
2
43749 43
0
9 Inverter~
13 1689 2581 0 2 22
0 55 3
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U21C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
999 0 0
2
43749 44
0
8 2-In OR~
219 1689 2533 0 3 22
0 56 39 55
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U20D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8787 0 0
2
43749 45
0
8 2-In OR~
219 1721 2456 0 3 22
0 5 21 56
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U20C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3348 0 0
2
43749 46
0
9 2-In AND~
219 1781 2366 0 3 22
0 40 38 5
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U24D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3395 0 0
2
43749 47
0
9 2-In AND~
219 1674 2344 0 3 22
0 40 44 21
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U24C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7740 0 0
2
43749 48
0
9 Inverter~
13 1489 2319 0 2 22
0 57 11
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U21B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
6480 0 0
2
43749 49
0
8 2-In OR~
219 1488 2273 0 3 22
0 39 8 57
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U20B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
342 0 0
2
43749 50
0
9 2-In AND~
219 1497 2197 0 3 22
0 58 45 39
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U24B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9953 0 0
2
43749 51
0
9 Inverter~
13 1353 2243 0 2 22
0 8 13
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U21A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
361 0 0
2
43749 52
0
9 Inverter~
13 1139 2264 0 2 22
0 59 10
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U18F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3343 0 0
2
43749 53
0
8 2-In OR~
219 1139 2177 0 3 22
0 54 7 59
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U20A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7923 0 0
2
43749 54
0
9 2-In AND~
219 1159 2108 0 3 22
0 45 40 54
0
0 0 608 270
5 74F08
-18 -24 17 -16
4 U19A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6174 0 0
2
43749 55
0
7 Ground~
168 588 1927 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6692 0 0
2
43749 56
0
7 74LS154
95 818 1901 0 22 45
0 2 2 61 62 63 60 107 108 109
110 111 112 113 114 115 116 46 47 48
49 50 51
0
0 0 4832 692
7 74LS154
-24 -87 25 -79
3 U15
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
8790 0 0
2
5.89911e-315 5.41378e-315
0
7 Ground~
168 1499 578 0 1 3
0 2
0
0 0 53344 692
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4595 0 0
2
43749 57
0
7 Ground~
168 1475 755 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
667 0 0
2
5.89911e-315 5.41896e-315
0
7 74LS157
122 1543 749 0 14 29
0 5 77 29 75 28 74 31 76 32
2 70 71 73 72
0
0 0 4320 270
7 74LS157
-24 -60 25 -52
3 U35
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8743 0 0
2
5.89911e-315 5.42414e-315
0
7 Ground~
168 1895 570 0 1 3
0 2
0
0 0 53344 180
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8298 0 0
2
5.89911e-315 5.42933e-315
0
7 74LS173
129 1836 642 0 14 29
0 2 2 2 27 66 67 68 65 2
2 76 74 75 77
0
0 0 4320 0
7 74LS173
-24 -51 25 -43
3 U34
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
313 0 0
2
5.89911e-315 5.43192e-315
0
14 Logic Display~
6 1013 1332 0 1 2
10 22
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L319
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7548 0 0
2
43749 58
0
14 Logic Display~
6 984 1332 0 1 2
10 23
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L318
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8973 0 0
2
43749 59
0
14 Logic Display~
6 954 1332 0 1 2
10 24
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L317
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9712 0 0
2
43749 60
0
14 Logic Display~
6 924 1332 0 1 2
10 25
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L316
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4518 0 0
2
43749 61
0
14 Logic Display~
6 867 1332 0 1 2
10 78
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L315
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5596 0 0
2
43749 62
0
14 Logic Display~
6 836 1332 0 1 2
10 79
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L314
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
692 0 0
2
43749 63
0
14 Logic Display~
6 804 1331 0 1 2
10 80
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L313
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6258 0 0
2
43749 64
0
14 Logic Display~
6 772 1331 0 1 2
10 81
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L312
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5578 0 0
2
43749 65
0
14 Logic Display~
6 772 962 0 1 2
10 81
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L311
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8709 0 0
2
43749 66
0
14 Logic Display~
6 804 962 0 1 2
10 80
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L310
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9131 0 0
2
43749 67
0
14 Logic Display~
6 836 962 0 1 2
10 79
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L309
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3645 0 0
2
43749 68
0
14 Logic Display~
6 867 962 0 1 2
10 78
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L308
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7613 0 0
2
43749 69
0
14 Logic Display~
6 924 962 0 1 2
10 25
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L307
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9467 0 0
2
43749 70
0
14 Logic Display~
6 954 962 0 1 2
10 24
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L306
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3932 0 0
2
43749 71
0
14 Logic Display~
6 984 962 0 1 2
10 23
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L305
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5288 0 0
2
43749 72
0
14 Logic Display~
6 1013 961 0 1 2
10 22
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L304
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4934 0 0
2
43749 73
0
14 Logic Display~
6 772 586 0 1 2
10 81
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L303
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5987 0 0
2
43749 74
0
14 Logic Display~
6 804 586 0 1 2
10 80
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L302
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7737 0 0
2
43749 75
0
14 Logic Display~
6 836 585 0 1 2
10 79
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L301
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4200 0 0
2
43749 76
0
14 Logic Display~
6 924 586 0 1 2
10 25
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L299
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5780 0 0
2
43749 77
0
14 Logic Display~
6 954 586 0 1 2
10 24
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L298
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6490 0 0
2
43749 78
0
14 Logic Display~
6 984 586 0 1 2
10 23
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L297
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8663 0 0
2
43749 79
0
14 Logic Display~
6 1013 586 0 1 2
10 22
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L296
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
318 0 0
2
43749 80
0
14 Logic Display~
6 612 274 0 1 2
10 22
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L287
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
348 0 0
2
43749 81
0
14 Logic Display~
6 612 256 0 1 2
10 23
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L286
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8551 0 0
2
43749 82
0
14 Logic Display~
6 612 238 0 1 2
10 24
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L285
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7295 0 0
2
43749 83
0
14 Logic Display~
6 612 220 0 1 2
10 25
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L284
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9900 0 0
2
43749 84
0
14 Logic Display~
6 488 274 0 1 2
10 83
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L283
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8725 0 0
2
43749 85
0
14 Logic Display~
6 488 256 0 1 2
10 84
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L282
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
366 0 0
2
43749 86
0
14 Logic Display~
6 488 238 0 1 2
10 85
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L281
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5762 0 0
2
43749 87
0
14 Logic Display~
6 488 220 0 1 2
10 86
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L280
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4943 0 0
2
43749 88
0
14 Logic Display~
6 722 345 0 1 2
10 22
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L275
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3435 0 0
2
43749 89
0
14 Logic Display~
6 700 327 0 1 2
10 23
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L274
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8705 0 0
2
43749 90
0
14 Logic Display~
6 673 308 0 1 2
10 24
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L273
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4331 0 0
2
43749 91
0
14 Logic Display~
6 649 292 0 1 2
10 25
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L272
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
787 0 0
2
43749 92
0
14 Logic Display~
6 608 635 0 1 2
10 87
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L263
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3655 0 0
2
43749 93
0
14 Logic Display~
6 590 635 0 1 2
10 88
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L262
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6682 0 0
2
43749 94
0
14 Logic Display~
6 572 635 0 1 2
10 89
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L261
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
582 0 0
2
43749 95
0
14 Logic Display~
6 554 635 0 1 2
10 90
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L260
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3125 0 0
2
43749 96
0
14 Logic Display~
6 745 707 0 1 2
10 22
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L259
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5466 0 0
2
43749 97
0
14 Logic Display~
6 745 698 0 1 2
10 23
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L258
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
52 0 0
2
43749 98
0
14 Logic Display~
6 745 689 0 1 2
10 24
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L257
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3898 0 0
2
43749 99
0
14 Logic Display~
6 745 680 0 1 2
10 25
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L256
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9413 0 0
2
43749 100
0
14 Logic Display~
6 745 671 0 1 2
10 78
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L255
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8576 0 0
2
43749 101
0
14 Logic Display~
6 745 662 0 1 2
10 79
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L254
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
622 0 0
2
43749 102
0
14 Logic Display~
6 745 653 0 1 2
10 80
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L253
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9152 0 0
2
43749 103
0
14 Logic Display~
6 745 644 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L252
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
783 0 0
2
43749 104
0
14 Logic Display~
6 705 1157 0 1 2
10 22
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L239
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4262 0 0
2
43749 105
0
14 Logic Display~
6 684 1148 0 1 2
10 23
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L238
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6121 0 0
2
43749 106
0
14 Logic Display~
6 665 1139 0 1 2
10 24
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L237
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3879 0 0
2
43749 107
0
14 Logic Display~
6 646 1130 0 1 2
10 25
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L236
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7345 0 0
2
43749 108
0
14 Logic Display~
6 471 1273 0 1 2
10 78
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L235
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3198 0 0
2
43749 109
0
14 Logic Display~
6 457 1263 0 1 2
10 79
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L234
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9849 0 0
2
43749 110
0
14 Logic Display~
6 446 1254 0 1 2
10 80
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L233
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
479 0 0
2
43749 111
0
14 Logic Display~
6 435 1244 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L232
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3905 0 0
2
43749 112
0
14 Logic Display~
6 510 1357 0 1 2
10 60
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L231
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4394 0 0
2
43749 113
0
14 Logic Display~
6 519 1336 0 1 2
10 63
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L230
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4391 0 0
2
43749 114
0
14 Logic Display~
6 528 1315 0 1 2
10 62
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L229
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3681 0 0
2
43749 115
0
14 Logic Display~
6 538 1299 0 1 2
10 61
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L228
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6466 0 0
2
43749 116
0
14 Logic Display~
6 757 1110 0 1 2
10 22
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L227
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5230 0 0
2
43749 117
0
14 Logic Display~
6 750 1101 0 1 2
10 23
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L226
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8324 0 0
2
43749 118
0
14 Logic Display~
6 739 1092 0 1 2
10 24
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L225
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3445 0 0
2
43749 119
0
14 Logic Display~
6 726 1083 0 1 2
10 25
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L224
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7543 0 0
2
43749 120
0
14 Logic Display~
6 1046 341 0 1 2
10 22
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L218
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
43749 121
0
14 Logic Display~
6 1046 323 0 1 2
10 23
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L217
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5476 0 0
2
43749 122
0
14 Logic Display~
6 1046 305 0 1 2
10 24
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L216
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3936 0 0
2
43749 123
0
14 Logic Display~
6 1046 287 0 1 2
10 25
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L215
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5770 0 0
2
43749 124
0
14 Logic Display~
6 1170 342 0 1 2
10 17
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L214
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7884 0 0
2
43749 125
0
14 Logic Display~
6 1170 323 0 1 2
10 14
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L213
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3690 0 0
2
43749 126
0
14 Logic Display~
6 1170 305 0 1 2
10 16
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L212
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3611 0 0
2
43749 127
0
14 Logic Display~
6 1169 287 0 1 2
10 15
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L211
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7912 0 0
2
43749 128
0
14 Logic Display~
6 1146 544 0 1 2
10 91
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L210
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6416 0 0
2
43749 129
0
14 Logic Display~
6 1146 526 0 1 2
10 92
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L209
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7278 0 0
2
43749 130
0
14 Logic Display~
6 1146 508 0 1 2
10 93
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L208
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6804 0 0
2
43749 131
0
14 Logic Display~
6 1146 490 0 1 2
10 94
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L207
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9568 0 0
2
43749 132
0
14 Logic Display~
6 1349 427 0 1 2
10 17
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L201
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7178 0 0
2
43749 133
0
14 Logic Display~
6 1335 427 0 1 2
10 14
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L200
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7982 0 0
2
43749 134
0
14 Logic Display~
6 1321 427 0 1 2
10 16
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L199
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
513 0 0
2
43749 135
0
14 Logic Display~
6 1308 427 0 1 2
10 15
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L198
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8190 0 0
2
43749 136
0
14 Logic Display~
6 1349 245 0 1 2
10 17
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L197
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5209 0 0
2
43749 137
0
14 Logic Display~
6 1335 245 0 1 2
10 14
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L196
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7239 0 0
2
43749 138
0
14 Logic Display~
6 1321 245 0 1 2
10 16
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L195
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9474 0 0
2
43749 139
0
14 Logic Display~
6 1308 245 0 1 2
10 15
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L194
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3783 0 0
2
43749 140
0
14 Logic Display~
6 1129 930 0 1 2
10 22
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L187
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5422 0 0
2
43749 141
0
14 Logic Display~
6 1108 921 0 1 2
10 23
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L186
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8527 0 0
2
43749 142
0
14 Logic Display~
6 1085 912 0 1 2
10 24
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L185
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
761 0 0
2
43749 143
0
14 Logic Display~
6 1065 902 0 1 2
10 25
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L184
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7323 0 0
2
43749 144
0
14 Logic Display~
6 1125 221 0 1 2
10 22
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L183
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8543 0 0
2
43749 145
0
14 Logic Display~
6 1101 212 0 1 2
10 23
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L182
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4240 0 0
2
43749 146
0
14 Logic Display~
6 1076 203 0 1 2
10 24
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L181
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7857 0 0
2
43749 147
0
14 Logic Display~
6 1055 194 0 1 2
10 25
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L180
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7255 0 0
2
43749 148
0
12 SPST Switch~
165 741 1470 0 10 11
0 95 27 0 0 0 0 0 0 0
1
0
0 0 4192 0
0
2 S7
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7736 0 0
2
43749 149
0
14 Logic Display~
6 2761 3065 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L174
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5435 0 0
2
5.89911e-315 5.43451e-315
0
14 Logic Display~
6 2732 2978 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L173
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3446 0 0
2
5.89911e-315 5.4371e-315
0
14 Logic Display~
6 2703 2902 0 1 2
10 117
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L172
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3914 0 0
2
5.89911e-315 5.43969e-315
0
14 Logic Display~
6 2671 2820 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L171
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3948 0 0
2
5.89911e-315 5.44228e-315
0
14 Logic Display~
6 2641 2746 0 1 2
10 118
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L170
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3901 0 0
2
5.89911e-315 5.44487e-315
0
14 Logic Display~
6 2611 2670 0 1 2
10 119
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L169
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
6295 0 0
2
5.89911e-315 5.44746e-315
0
14 Logic Display~
6 2581 2598 0 1 2
10 120
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L168
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
332 0 0
2
5.89911e-315 5.45005e-315
0
14 Logic Display~
6 2551 2530 0 1 2
10 121
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L167
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
9737 0 0
2
5.89911e-315 5.45264e-315
0
14 Logic Display~
6 2522 2448 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L166
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9910 0 0
2
5.89911e-315 5.45523e-315
0
14 Logic Display~
6 2463 2290 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L164
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
2
5.89911e-315 5.45782e-315
0
14 Logic Display~
6 2762 2258 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L163
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3138 0 0
2
5.89911e-315 5.46041e-315
0
14 Logic Display~
6 2731 2236 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L162
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5409 0 0
2
5.89911e-315 5.463e-315
0
14 Logic Display~
6 2704 2214 0 1 2
10 122
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L161
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
983 0 0
2
5.89911e-315 5.46559e-315
0
14 Logic Display~
6 2671 2188 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L160
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6652 0 0
2
5.89911e-315 5.46818e-315
0
14 Logic Display~
6 2522 2074 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L155
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4281 0 0
2
5.89911e-315 5.47077e-315
0
14 Logic Display~
6 2463 2018 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L153
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6847 0 0
2
5.89911e-315 5.47207e-315
0
14 Logic Display~
6 2761 1730 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L152
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6543 0 0
2
5.89911e-315 5.47336e-315
0
14 Logic Display~
6 2732 1714 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L151
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89911e-315 5.47466e-315
0
14 Logic Display~
6 2670 1678 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L149
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3828 0 0
2
5.89911e-315 5.47595e-315
0
14 Logic Display~
6 2522 1598 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L144
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
955 0 0
2
5.89911e-315 5.47725e-315
0
14 Logic Display~
6 2463 1531 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L142
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7782 0 0
2
5.89911e-315 5.47854e-315
0
14 Logic Display~
6 2463 1531 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L141
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
824 0 0
2
5.89911e-315 5.47984e-315
0
14 Logic Display~
6 2762 1307 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L140
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6983 0 0
2
5.89911e-315 5.48113e-315
0
14 Logic Display~
6 2733 1286 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L139
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3185 0 0
2
5.89911e-315 5.48243e-315
0
14 Logic Display~
6 2671 1251 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L137
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4213 0 0
2
5.89911e-315 5.48372e-315
0
14 Logic Display~
6 2522 1152 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L132
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9765 0 0
2
5.89911e-315 5.48502e-315
0
14 Logic Display~
6 2463 1113 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L130
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8986 0 0
2
5.89911e-315 5.48631e-315
0
14 Logic Display~
6 2761 544 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L129
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3273 0 0
2
5.89911e-315 5.48761e-315
0
14 Logic Display~
6 2732 520 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L128
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5636 0 0
2
5.89911e-315 5.4889e-315
0
14 Logic Display~
6 2671 470 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L126
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
327 0 0
2
5.89911e-315 5.4902e-315
0
14 Logic Display~
6 2522 505 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L121
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9233 0 0
2
5.89911e-315 5.49149e-315
0
14 Logic Display~
6 2761 903 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L120
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3875 0 0
2
5.89911e-315 5.49279e-315
0
14 Logic Display~
6 2732 882 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L119
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9991 0 0
2
5.89911e-315 5.49408e-315
0
14 Logic Display~
6 2671 847 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L117
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
5.89911e-315 5.49538e-315
0
14 Logic Display~
6 2522 732 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L112
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8874 0 0
2
5.89911e-315 5.49667e-315
0
14 Logic Display~
6 27 2738 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L110
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7400 0 0
2
5.89911e-315 5.49797e-315
0
14 Logic Display~
6 57 2680 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L109
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3623 0 0
2
5.89911e-315 5.49926e-315
0
14 Logic Display~
6 85 2616 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L108
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3311 0 0
2
5.89911e-315 5.50056e-315
0
14 Logic Display~
6 113 2552 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L107
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5736 0 0
2
5.89911e-315 5.50185e-315
0
14 Logic Display~
6 169 2424 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L105
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3143 0 0
2
5.89911e-315 5.50315e-315
0
14 Logic Display~
6 196 2363 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L104
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5835 0 0
2
5.89911e-315 5.50444e-315
0
14 Logic Display~
6 223 2309 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L103
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5108 0 0
2
5.89911e-315 5.50574e-315
0
14 Logic Display~
6 224 2044 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L102
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3320 0 0
2
5.89911e-315 5.50703e-315
0
14 Logic Display~
6 196 1997 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L101
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.89911e-315 5.50833e-315
0
14 Logic Display~
6 169 1949 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L100
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3557 0 0
2
5.89911e-315 5.50963e-315
0
14 Logic Display~
6 113 1832 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L98
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7246 0 0
2
5.89911e-315 5.51092e-315
0
14 Logic Display~
6 86 1776 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L97
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3916 0 0
2
5.89911e-315 5.51222e-315
0
14 Logic Display~
6 57 1726 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L96
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
614 0 0
2
5.89911e-315 5.51286e-315
0
14 Logic Display~
6 28 1686 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L95
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8494 0 0
2
5.89911e-315 5.51351e-315
0
14 Logic Display~
6 223 1432 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L94
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
774 0 0
2
5.89911e-315 5.51416e-315
0
14 Logic Display~
6 196 1376 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L93
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
715 0 0
2
5.89911e-315 5.51481e-315
0
14 Logic Display~
6 169 1330 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L92
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3281 0 0
2
5.89911e-315 5.51545e-315
0
14 Logic Display~
6 115 1248 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L90
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
5.89911e-315 5.5161e-315
0
14 Logic Display~
6 85 1212 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L89
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7233 0 0
2
5.89911e-315 5.51675e-315
0
14 Logic Display~
6 57 1166 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L88
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3410 0 0
2
5.89911e-315 5.5174e-315
0
14 Logic Display~
6 28 1122 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L87
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3616 0 0
2
5.89911e-315 5.51804e-315
0
14 Logic Display~
6 223 1173 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L86
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5202 0 0
2
5.89911e-315 5.51869e-315
0
14 Logic Display~
6 196 1008 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L85
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9145 0 0
2
5.89911e-315 5.51934e-315
0
14 Logic Display~
6 169 906 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L84
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9815 0 0
2
5.89911e-315 5.51999e-315
0
14 Logic Display~
6 114 824 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L82
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4766 0 0
2
5.89911e-315 5.52063e-315
0
14 Logic Display~
6 86 770 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L81
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8325 0 0
2
5.89911e-315 5.52128e-315
0
14 Logic Display~
6 57 731 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L80
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7196 0 0
2
5.89911e-315 5.52193e-315
0
14 Logic Display~
6 28 707 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L79
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3567 0 0
2
5.89911e-315 5.52258e-315
0
14 Logic Display~
6 532 105 0 1 2
10 7
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L74
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5877 0 0
2
5.89911e-315 5.52517e-315
0
14 Logic Display~
6 194 104 0 1 2
10 7
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L73
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4785 0 0
2
5.89911e-315 5.52581e-315
0
14 Logic Display~
6 159 206 0 1 2
10 8
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L72
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3822 0 0
2
5.89911e-315 5.52646e-315
0
14 Logic Display~
6 193 301 0 1 2
10 10
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L70
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7640 0 0
2
5.89911e-315 5.52711e-315
0
14 Logic Display~
6 189 641 0 1 2
10 34
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L69
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9221 0 0
2
5.89911e-315 5.52776e-315
0
14 Logic Display~
6 189 670 0 1 2
10 11
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L68
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6484 0 0
2
5.89911e-315 5.52841e-315
0
14 Logic Display~
6 1729 473 0 1 2
10 2
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L65
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3689 0 0
2
5.89911e-315 5.5297e-315
0
14 Logic Display~
6 1692 464 0 1 2
10 18
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L64
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3952 0 0
2
5.89911e-315 5.53035e-315
0
14 Logic Display~
6 1650 455 0 1 2
10 123
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L63
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3631 0 0
2
5.89911e-315 5.531e-315
0
14 Logic Display~
6 1610 445 0 1 2
10 2
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L62
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9359 0 0
2
5.89911e-315 5.53164e-315
0
14 Logic Display~
6 1607 266 0 1 2
10 4
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L58
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5584 0 0
2
5.89911e-315 5.53423e-315
0
9 Terminal~
194 2761 3121 0 1 3
0 3
0
0 0 49504 180
5 LaBAR
6 -7 41 1
3 T19
-11 -32 10 -24
0
6 LaBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4973 0 0
2
43749 150
0
9 Terminal~
194 2732 3039 0 1 3
0 4
0
0 0 49504 180
2 Ea
-5 -1 9 7
3 T18
-10 -32 11 -24
0
3 Ea;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3239 0 0
2
43749 151
0
9 Terminal~
194 2704 2956 0 1 3
0 0
0
0 0 49504 180
2 Eu
-5 1 9 9
3 T17
-10 -32 11 -24
0
3 Eu;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
4244 0 0
2
43749 152
0
9 Terminal~
194 2671 2872 0 1 3
0 5
0
0 0 49504 180
1 M
-3 -1 4 7
3 T16
-11 -32 10 -24
0
2 M;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3391 0 0
2
43749 153
0
9 Terminal~
194 2641 2800 0 1 3
0 0
0
0 0 49504 180
3 Cin
-9 -1 12 7
3 T15
-11 -32 10 -24
0
4 Cin;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
4243 0 0
2
43749 154
0
9 Terminal~
194 2611 2731 0 1 3
0 0
0
0 0 49504 180
2 S3
-6 -2 8 6
3 T14
-10 -32 11 -24
0
3 S3;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
3907 0 0
2
43749 155
0
9 Terminal~
194 2582 2652 0 1 3
0 0
0
0 0 49504 180
2 S2
-5 0 9 8
3 T13
-10 -32 11 -24
0
3 S2;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
728 0 0
2
43749 156
0
9 Terminal~
194 2576 2776 0 1 3
0 0
0
0 0 49504 180
2 S1
-6 -1 8 7
3 T12
-10 -32 11 -24
0
3 S1;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
3585 0 0
2
43749 157
0
9 Terminal~
194 2522 2497 0 1 3
0 5
0
0 0 49504 180
2 S0
7 -7 21 1
3 T11
-10 -32 11 -24
0
3 S0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3565 0 0
2
43749 158
0
9 Terminal~
194 2464 2337 0 1 3
0 6
0
0 0 49504 692
5 LoBAR
-16 -1 19 7
2 T9
-8 -32 6 -24
0
6 LoBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3966 0 0
2
43749 159
0
9 Terminal~
194 28 2783 0 1 3
0 7
0
0 0 49504 180
2 Ep
-7 0 7 8
2 T8
-7 -32 7 -24
0
3 Ep;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3714 0 0
2
43749 160
0
9 Terminal~
194 57 2720 0 1 3
0 8
0
0 0 49504 180
2 Cp
-6 0 8 8
2 T7
-7 -32 7 -24
0
3 Cp;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3406 0 0
2
43749 161
0
9 Terminal~
194 86 2662 0 1 3
0 9
0
0 0 49504 180
5 LpBAR
-16 -1 19 7
2 T6
-7 -32 7 -24
0
6 LpBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3132 0 0
2
43749 162
0
9 Terminal~
194 114 2600 0 1 3
0 10
0
0 0 49504 180
5 LmBAR
-16 -1 19 7
2 T5
-8 -32 6 -24
0
6 LmBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3842 0 0
2
43749 163
0
9 Terminal~
194 169 2470 0 1 3
0 11
0
0 0 49504 180
5 CEbar
-17 -1 18 7
2 T3
-8 -32 6 -24
0
6 CEbar;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6183 0 0
2
43749 164
0
9 Terminal~
194 226 2473 0 1 3
0 12
0
0 0 49504 180
5 EiBAR
-16 -1 19 7
2 T2
-8 -32 6 -24
0
6 EiBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3356 0 0
2
43749 165
0
9 Terminal~
194 223 2354 0 1 3
0 13
0
0 0 49504 180
5 LiBAR
-17 -1 18 7
2 T1
-7 -32 7 -24
0
6 LiBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3525 0 0
2
43749 166
0
14 Logic Display~
6 927 1623 0 1 2
10 7
0
0 0 53360 270
6 100MEG
3 -16 45 -8
3 L10
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
43749 167
0
14 Logic Display~
6 927 1650 0 1 2
10 8
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L9
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
346 0 0
2
43749 168
0
14 Logic Display~
6 927 1680 0 1 2
10 40
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L8
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3169 0 0
2
43749 169
0
14 Logic Display~
6 927 1708 0 1 2
10 58
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L7
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4826 0 0
2
43749 170
0
14 Logic Display~
6 2288 1709 0 1 2
10 58
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L14
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3971 0 0
2
5.89911e-315 5.53488e-315
0
14 Logic Display~
6 2287 1681 0 1 2
10 40
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L13
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3607 0 0
2
5.89911e-315 5.53553e-315
0
14 Logic Display~
6 2287 1651 0 1 2
10 8
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L12
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3506 0 0
2
5.89911e-315 5.53618e-315
0
14 Logic Display~
6 2287 1624 0 1 2
10 7
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L11
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7829 0 0
2
5.89911e-315 5.53682e-315
0
14 Logic Display~
6 1025 1434 0 1 2
10 95
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3890 0 0
2
43749 171
0
7 74LS107
112 1439 1476 0 12 25
0 100 58 95 97 7 99 95 97 99
7 8 98
0
0 0 4320 0
7 74LS107
-24 -51 25 -43
3 U17
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 4 12 13 8 11 9 10 3
2 5 6 1 4 12 13 8 11 9
10 3 2 5 6 0
65 0 0 0 1 1 0 0
1 U
3126 0 0
2
43749 172
0
7 74LS107
112 1214 1479 0 12 25
0 8 98 95 97 40 101 95 97 40
101 58 100
0
0 0 4320 0
7 74LS107
-24 -51 25 -43
3 U16
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 4 12 13 8 11 9 10 3
2 5 6 1 4 12 13 8 11 9
10 3 2 5 6 0
65 0 0 0 1 0 0 0
1 U
3935 0 0
2
43749 173
0
14 Logic Display~
6 221 32 0 1 2
10 27
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9746 0 0
2
43749 174
0
7 Pulser~
4 158 73 0 11 12
0 35 124 27 125 0 0 10 10 -1
7 1
0
0 0 4128 0
0
3 V11
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7330 0 0
2
43749 175
0
7 74LS126
116 558 241 0 12 25
0 7 86 7 85 7 84 7 83 25
24 23 22
0
0 0 4832 0
7 74LS126
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3972 0 0
2
43749 176
0
7 74LS193
137 393 227 0 14 29
0 27 8 9 102 25 24 23 22 126
127 86 85 84 83
0
0 0 4320 0
7 74LS193
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7818 0 0
2
43749 177
0
7 74LS173
129 598 354 0 14 29
0 2 10 10 27 25 24 23 22 2
2 90 89 88 87
0
0 0 4320 782
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3818 0 0
2
43749 178
0
7 74LS173
129 1253 188 0 14 29
0 2 3 3 27 25 24 23 22 2
2 15 16 14 17
0
0 0 4320 0
7 74LS173
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
8835 0 0
2
43749 179
0
7 74LS126
116 1103 309 0 12 25
0 4 15 4 16 4 14 4 17 25
24 23 22
0
0 0 4320 512
7 74LS126
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
7484 0 0
2
43749 180
0
7 74LS126
116 1105 512 0 12 25
0 20 94 20 93 20 92 20 91 25
24 23 22
0
0 0 4320 512
7 74LS126
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
792 0 0
2
43749 181
0
7 74LS181
132 1249 494 0 22 45
0 2 19 18 2 15 16 14 17 72
73 71 70 96 5 128 129 130 131 94
93 92 91
0
0 0 12512 512
7 74LS181
-24 -69 25 -61
2 U7
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 254
65 0 0 512 1 0 0 0
1 U
3826 0 0
2
43749 182
0
7 74LS173
129 1272 713 0 14 29
0 2 33 33 27 25 24 23 22 2
2 32 31 28 29
0
0 0 4320 0
7 74LS173
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7958 0 0
2
43749 183
0
7 Ground~
168 534 322 0 1 3
0 2
0
0 0 53344 270
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6736 0 0
2
43749 184
0
7 Ground~
168 1305 169 0 1 3
0 2
0
0 0 53344 782
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3755 0 0
2
43749 185
0
7 Ground~
168 1284 605 0 1 3
0 2
0
0 0 53344 692
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
397 0 0
2
43749 186
0
6 1K RAM
79 658 666 0 20 41
0 82 82 82 82 82 82 90 89 88
87 81 80 79 78 25 24 23 22 11
34
0
0 0 4320 0
5 RAM1K
-17 -19 18 -11
3 U11
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 1 0 0 0
1 U
5190 0 0
2
43749 187
0
7 74LS173
129 471 1191 0 14 29
0 2 13 13 27 81 80 79 78 2
2 61 62 63 60
0
0 0 4320 0
7 74LS173
-24 -51 25 -43
3 U13
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
9188 0 0
2
43749 188
0
7 Ground~
168 526 1163 0 1 3
0 2
0
0 0 53344 782
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3651 0 0
2
43749 189
0
7 Ground~
168 627 1036 0 1 3
0 2
0
0 0 53344 692
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3415 0 0
2
43749 190
0
7 74LS173
129 675 1077 0 14 29
0 2 13 13 27 25 24 23 22 12
12 25 24 23 22
0
0 0 4320 0
7 74LS173
-24 -51 25 -43
3 U14
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7597 0 0
2
43749 191
0
14 Logic Display~
6 1420 878 0 1 2
10 104
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
350 0 0
2
43749 192
0
14 Logic Display~
6 1443 878 0 1 2
10 103
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3153 0 0
2
43749 193
0
14 Logic Display~
6 1397 878 0 1 2
10 105
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
634 0 0
2
43749 194
0
14 Logic Display~
6 1374 878 0 1 2
10 106
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8956 0 0
2
43749 195
0
7 Ground~
168 1293 838 0 1 3
0 2
0
0 0 53344 692
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3342 0 0
2
43749 196
0
7 74LS173
129 1255 897 0 14 29
0 2 6 6 27 25 24 23 22 2
2 106 105 104 103
0
0 0 4320 0
7 74LS173
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
2
43749 197
0
601
1 0 14 0 0 0 0 14 0 0 5 2
1598 187
1598 187
1 0 15 0 0 0 0 16 0 0 3 2
1531 184
1531 184
0 0 15 0 0 4224 0 0 0 582 0 3
1308 199
1531 199
1531 178
0 1 16 0 0 4224 0 0 15 581 0 3
1321 209
1567 209
1567 186
0 0 14 0 0 4224 0 0 0 580 0 3
1335 216
1598 216
1598 184
0 1 17 0 0 4224 0 0 13 579 0 4
1349 226
1626 226
1626 184
1625 184
0 0 5 0 0 4096 0 0 0 484 257 2
1709 381
1919 381
1 0 18 0 0 4096 0 2 0 0 252 2
1886 498
1886 499
2 1 19 0 0 4224 0 282 3 0 0 3
1281 458
1912 458
1912 457
0 0 20 0 0 8192 0 0 0 11 0 3
2701 360
2701 361
2317 361
0 0 20 0 0 4224 0 0 0 12 0 2
2701 1667
2701 350
3 0 20 0 0 0 0 17 0 0 0 4
2274 2633
2274 2722
2701 2722
2701 1663
0 2 5 0 0 0 0 0 17 97 0 4
2337 2536
2266 2536
2266 2587
2265 2587
0 1 21 0 0 4224 0 0 17 120 0 4
1672 2410
2300 2410
2300 2587
2283 2587
1 0 2 0 0 0 0 19 0 0 27 2
1789 492
1789 492
0 12 22 0 0 12288 0 0 281 595 0 6
1013 548
1019 548
1019 563
1068 563
1068 548
1073 548
0 11 23 0 0 4096 0 0 281 594 0 2
984 530
1073 530
0 10 24 0 0 4096 0 0 281 490 0 2
1000 512
1073 512
0 9 25 0 0 8192 0 0 281 0 0 3
1059 496
1059 494
1073 494
0 0 26 0 0 4224 0 0 0 0 0 4
2406 612
2417 612
2417 613
2418 613
0 0 27 0 0 4096 27 0 0 247 217 2
357 67
599 67
0 0 25 0 0 4096 0 0 0 178 597 2
1078 642
924 642
0 0 24 0 0 4096 0 0 0 179 596 2
1084 731
954 731
0 0 23 0 0 4096 0 0 0 180 594 2
1090 761
984 761
0 0 22 0 0 4096 0 0 0 181 595 2
1087 791
1013 791
1 0 2 0 0 0 0 241 0 0 27 2
1744 476
1744 476
4 0 2 0 0 4096 0 282 0 0 0 5
1281 476
1769 476
1769 492
1796 492
1796 496
1 0 28 0 0 0 0 20 0 0 30 2
1469 661
1469 661
1 0 29 0 0 0 0 21 0 0 204 2
1467 690
1467 690
13 5 28 0 0 4224 0 283 77 0 0 5
1304 740
1439 740
1439 661
1542 661
1542 722
0 0 30 0 0 4224 0 0 0 0 0 4
1304 740
1439 740
1439 661
1445 661
1 0 2 0 0 0 0 75 0 0 174 2
1499 586
1500 589
1 0 31 0 0 4096 0 22 0 0 203 2
1436 639
1436 641
1 0 32 0 0 4096 0 23 0 0 202 2
1435 602
1435 601
1 0 33 0 0 4096 0 24 0 0 36 2
1530 519
1530 517
0 0 33 0 0 41088 0 0 0 565 104 12
1217 650
1184 650
1184 581
1464 581
1464 517
1769 517
1769 539
2220 539
2220 570
2874 570
2874 2660
1967 2660
2 0 6 0 0 8192 0 25 0 0 482 3
2357 2200
2357 2202
2464 2202
0 0 34 0 0 4096 0 0 0 161 262 2
143 693
143 713
2 0 9 0 0 16384 0 26 0 0 0 5
2539 2693
2539 2692
2546 2692
2546 2903
2004 2903
1 0 35 0 0 8320 0 275 0 0 165 3
134 64
134 67
110 67
0 0 27 0 0 0 27 0 0 164 486 2
278 242
278 357
0 1 36 0 0 4224 0 0 25 100 0 3
2092 2202
2321 2202
2321 2200
0 0 3 0 0 12288 0 0 0 116 481 8
1692 2642
1750 2642
1750 3040
2535 3040
2535 3056
2739 3056
2739 3050
2761 3050
0 0 4 0 0 8192 0 0 0 99 259 7
2133 2664
2133 2994
2635 2994
2635 3027
2670 3027
2670 3013
2732 3013
0 0 12 0 0 4096 0 0 0 108 46 3
1837 2667
1026 2667
1026 2465
0 0 12 0 0 0 0 0 0 261 0 4
226 2428
580 2428
580 2465
1038 2465
0 0 9 0 0 4096 0 0 0 48 480 6
1115 2903
79 2903
79 2764
93 2764
93 2471
86 2471
0 0 9 0 0 0 0 0 0 39 0 2
2007 2903
1110 2903
0 1 37 0 0 4096 0 0 26 62 0 3
2482 2692
2503 2692
2503 2693
0 0 9 0 0 0 0 0 0 480 175 5
86 735
86 357
96 357
96 218
349 218
0 0 5 0 0 4096 0 0 0 97 257 2
2337 2484
2671 2484
0 0 5 0 0 0 0 0 0 97 483 2
2337 2403
2522 2403
0 0 11 0 0 4096 0 0 0 54 253 2
543 2268
169 2268
0 0 11 0 0 4096 0 0 0 128 0 4
1492 2376
618 2376
618 2268
540 2268
0 0 13 0 0 4096 0 0 0 136 260 4
1356 2346
642 2346
642 2238
223 2238
0 0 8 0 0 12288 0 0 0 139 479 4
1260 2325
682 2325
682 2211
57 2211
0 0 10 0 0 8192 0 0 0 58 254 3
740 2305
740 2179
114 2179
0 0 10 0 0 0 0 0 0 141 0 2
1142 2305
737 2305
0 0 7 0 0 4096 0 0 0 151 255 2
1100 2090
28 2090
2 0 38 0 0 12288 0 64 0 0 76 4
1770 2344
1770 2339
1733 2339
1733 1861
0 2 39 0 0 4224 0 0 62 127 0 4
1602 2243
1602 2468
1683 2468
1683 2517
0 1 37 0 0 8192 0 0 39 63 0 5
2434 2580
2482 2580
2482 2694
2489 2694
2489 2704
0 1 37 0 0 4224 0 0 42 111 0 5
1919 2434
2434 2434
2434 2637
2431 2637
2431 2677
0 0 40 0 0 4096 0 0 0 114 115 3
1899 2340
1899 2282
1881 2282
0 1 41 0 0 4096 0 0 55 74 0 4
2107 1949
2107 2128
2101 2128
2101 2138
2 0 42 0 0 4096 0 58 0 0 77 2
2054 2456
2054 1836
1 0 43 0 0 4096 0 60 0 0 75 2
1917 2371
1917 1905
1 0 41 0 0 0 0 27 0 0 74 2
1039 1949
1039 1949
1 0 43 0 0 0 0 28 0 0 75 2
1037 1905
1037 1905
1 0 38 0 0 0 0 29 0 0 76 2
1036 1862
1036 1861
1 0 42 0 0 0 0 30 0 0 77 2
1036 1837
1036 1836
1 0 44 0 0 4096 0 31 0 0 78 2
1034 1806
1034 1805
1 0 45 0 0 4096 0 32 0 0 79 2
1024 1776
1024 1775
2 0 41 0 0 4224 0 33 0 0 0 2
1012 1949
2369 1949
2 0 43 0 0 4224 0 34 0 0 0 2
1013 1905
2364 1905
2 0 38 0 0 4224 0 35 0 0 0 2
1023 1861
2383 1861
2 0 42 0 0 4224 0 36 0 0 0 2
1022 1836
2378 1836
2 0 44 0 0 4224 0 37 0 0 0 2
983 1805
2376 1805
2 0 45 0 0 4224 0 38 0 0 0 2
979 1775
2371 1775
17 1 46 0 0 4224 0 74 33 0 0 4
856 1878
927 1878
927 1949
976 1949
18 1 47 0 0 4224 0 74 34 0 0 5
856 1869
945 1869
945 1903
977 1903
977 1905
19 1 48 0 0 4224 0 74 35 0 0 3
856 1860
987 1860
987 1861
20 1 49 0 0 4224 0 74 36 0 0 4
856 1851
958 1851
958 1836
986 1836
21 1 50 0 0 4224 0 74 37 0 0 5
856 1842
917 1842
917 1804
947 1804
947 1805
22 1 51 0 0 8320 0 74 38 0 0 4
856 1833
891 1833
891 1775
943 1775
1 0 5 0 0 0 0 41 0 0 96 2
2372 2672
2370 2672
1 0 5 0 0 0 0 43 0 0 97 2
2338 2674
2337 2674
1 0 33 0 0 0 0 46 0 0 104 2
1968 2684
1967 2684
1 0 12 0 0 0 0 47 0 0 108 2
1838 2682
1837 2682
1 0 11 0 0 0 0 49 0 0 128 2
1494 2692
1492 2692
1 0 13 0 0 0 0 50 0 0 94 2
1358 2708
1356 2708
1 0 8 0 0 0 0 51 0 0 139 3
1259 2562
1260 2562
1260 2732
1 0 10 0 0 0 0 52 0 0 141 3
1163 2494
1163 2722
1141 2722
0 0 13 0 0 0 0 0 0 136 0 2
1356 2397
1356 2716
0 1 5 0 0 0 0 0 40 96 0 4
2370 2606
2396 2606
2396 2677
2398 2677
0 0 5 0 0 0 0 0 0 97 0 3
2337 2601
2370 2601
2370 2677
0 0 5 0 0 4096 0 0 0 121 0 3
1779 2399
2337 2399
2337 2680
0 1 36 0 0 0 0 0 44 100 0 6
2152 2490
2204 2490
2204 2653
2159 2653
2159 2681
2158 2681
3 1 4 0 0 0 0 54 45 0 0 5
2143 2573
2143 2664
2071 2664
2071 2686
2072 2686
3 1 36 0 0 0 0 55 54 0 0 6
2092 2183
2092 2286
2154 2286
2154 2483
2152 2483
2152 2527
0 2 52 0 0 4224 0 0 54 105 0 3
2064 2510
2134 2510
2134 2527
2 0 40 0 0 0 0 55 0 0 103 3
2083 2138
2084 2138
2084 2098
0 0 40 0 0 4096 0 0 0 448 0 2
2084 1684
2084 2103
2 0 33 0 0 0 0 56 0 0 0 4
2064 2571
2064 2623
1967 2623
1967 2689
1 3 52 0 0 0 0 56 58 0 0 3
2064 2535
2064 2501
2063 2501
1 3 53 0 0 8320 0 57 59 0 0 3
1924 2528
1924 2527
1926 2527
0 1 40 0 0 4096 0 0 58 448 0 5
2030 1684
2030 2307
2087 2307
2087 2456
2072 2456
0 0 12 0 0 0 0 0 0 109 0 2
1837 2603
1837 2687
2 0 12 0 0 0 0 57 0 0 0 3
1924 2564
1924 2603
1826 2603
0 0 54 0 0 4096 0 0 0 0 113 2
1949 2143
1949 2140
3 2 37 0 0 0 0 60 59 0 0 4
1908 2416
1919 2416
1919 2481
1917 2481
0 1 54 0 0 4096 0 0 59 113 0 3
1946 2140
1946 2481
1935 2481
0 0 54 0 0 4224 0 0 0 146 0 2
1151 2140
2010 2140
0 2 40 0 0 0 0 0 60 0 0 2
1899 2334
1899 2371
0 0 40 0 0 0 0 0 0 448 0 4
1853 1684
1853 2087
1881 2087
1881 2339
2 1 3 0 0 0 0 61 48 0 0 3
1692 2599
1692 2678
1690 2678
1 3 55 0 0 0 0 61 62 0 0 2
1692 2563
1692 2563
3 1 56 0 0 8320 0 63 62 0 0 4
1724 2486
1724 2506
1701 2506
1701 2517
2 0 21 0 0 0 0 63 0 0 120 2
1715 2440
1714 2440
3 0 21 0 0 0 0 65 0 0 0 4
1672 2367
1672 2420
1714 2420
1714 2444
3 1 5 0 0 0 0 64 63 0 0 4
1779 2389
1779 2416
1733 2416
1733 2440
1 0 40 0 0 0 0 64 0 0 123 2
1788 2344
1790 2344
0 0 40 0 0 0 0 0 0 124 0 7
1699 2237
1836 2237
1836 2307
1771 2307
1771 2333
1790 2333
1790 2349
0 1 40 0 0 0 0 0 65 448 0 4
1699 1684
1699 2283
1681 2283
1681 2322
2 0 44 0 0 0 0 65 0 0 126 2
1663 2322
1664 2322
0 0 44 0 0 0 0 0 0 78 0 2
1664 1805
1664 2330
0 0 39 0 0 0 0 0 0 132 0 2
1500 2243
1640 2243
2 0 11 0 0 0 0 66 0 0 0 2
1492 2337
1492 2696
1 3 57 0 0 4224 0 66 67 0 0 3
1492 2301
1492 2303
1491 2303
0 0 8 0 0 0 0 0 0 135 131 3
1443 2104
1469 2104
1469 2117
0 2 8 0 0 0 0 0 67 0 0 4
1469 2111
1469 2224
1482 2224
1482 2257
3 1 39 0 0 0 0 68 67 0 0 4
1495 2220
1495 2235
1500 2235
1500 2257
0 1 58 0 0 4096 0 0 68 462 0 3
1519 1712
1519 2175
1504 2175
0 2 45 0 0 0 0 0 68 79 0 3
1487 1775
1487 2175
1486 2175
0 0 8 0 0 0 0 0 0 139 0 2
1260 2104
1466 2104
2 0 13 0 0 0 0 69 0 0 0 2
1356 2261
1356 2401
1 0 8 0 0 0 0 69 0 0 138 2
1356 2225
1356 2225
0 0 8 0 0 0 0 0 0 139 0 3
1260 2146
1356 2146
1356 2229
0 0 8 0 0 4096 0 0 0 463 0 2
1260 1654
1260 2736
0 0 8 0 0 0 0 0 0 463 463 2
1188 1654
1241 1654
2 0 10 0 0 0 0 70 0 0 0 4
1142 2282
1142 2716
1141 2716
1141 2726
1 0 59 0 0 0 0 70 0 0 143 2
1142 2246
1142 2246
3 0 59 0 0 4224 0 71 0 0 0 2
1142 2207
1142 2250
0 1 7 0 0 0 0 0 53 151 0 3
1100 2164
1100 2733
1099 2733
0 2 7 0 0 0 0 0 71 151 0 3
1100 2036
1133 2036
1133 2161
1 3 54 0 0 0 0 71 72 0 0 4
1151 2161
1151 2140
1157 2140
1157 2131
2 0 40 0 0 0 0 72 0 0 150 2
1148 2086
1149 2086
1 0 45 0 0 0 0 72 0 0 149 2
1166 2086
1164 2086
0 0 45 0 0 0 0 0 0 79 0 2
1164 1775
1164 2091
0 0 40 0 0 0 0 0 0 448 0 2
1149 1684
1149 2091
0 0 7 0 0 0 0 0 0 464 0 2
1100 1627
1100 2172
1 0 2 0 0 0 0 73 0 0 153 2
588 1921
588 1923
0 0 2 0 0 0 0 0 0 154 0 2
726 1923
583 1923
1 2 2 0 0 0 0 74 74 0 0 4
780 1923
721 1923
721 1914
780 1914
0 0 60 0 0 4096 0 0 0 160 0 2
570 1860
539 1860
0 0 61 0 0 4096 0 0 0 0 157 4
469 1892
525 1892
525 1887
550 1887
3 0 61 0 0 4096 0 74 0 0 0 2
786 1887
544 1887
4 0 62 0 0 4096 0 74 0 0 0 4
786 1878
508 1878
508 1881
493 1881
5 0 63 0 0 4096 0 74 0 0 0 4
786 1869
540 1869
540 1871
513 1871
6 0 60 0 0 4096 0 74 0 0 0 2
786 1860
539 1860
0 20 34 0 0 16512 0 0 287 0 0 9
143 701
143 662
141 662
141 644
501 644
501 591
708 591
708 639
696 639
0 3 3 0 0 0 0 0 279 481 0 4
1867 108
1167 108
1167 179
1215 179
0 4 27 0 0 4096 27 0 79 488 0 4
1417 617
1750 617
1750 642
1804 642
0 0 27 0 0 0 27 0 0 0 247 2
278 257
278 200
1 0 35 0 0 0 0 12 0 0 0 2
101 67
114 67
0 1 35 0 0 0 0 0 12 0 0 2
106 67
101 67
0 0 64 0 0 4224 0 0 0 0 0 3
1887 452
1882 452
1882 456
1 1 2 0 0 16512 0 18 282 0 0 5
1883 416
1883 417
1856 417
1856 449
1281 449
0 1 5 0 0 4096 0 0 77 483 0 3
2522 689
1578 689
1578 722
0 0 58 0 0 0 0 0 0 462 462 2
1269 1712
1273 1712
0 2 8 0 0 0 0 0 277 263 0 4
69 239
69 208
361 208
361 209
0 0 12 0 0 0 0 0 0 0 261 5
196 1106
196 1091
180 1091
180 1204
196 1204
0 0 11 0 0 0 0 0 0 0 248 3
177 748
168 748
168 735
0 0 2 0 0 0 0 0 0 192 0 7
1782 632
1764 632
1764 564
1642 564
1642 589
1500 589
1500 584
3 0 9 0 0 0 0 277 0 0 0 2
355 218
345 218
0 0 62 0 0 0 0 0 0 471 158 4
528 1662
528 1787
745 1787
745 1878
1 8 65 0 0 12416 0 4 79 0 0 5
1803 1001
1803 1002
1790 1002
1790 678
1804 678
5 0 25 0 0 0 0 283 0 0 0 6
1240 722
1157 722
1157 642
1076 642
1076 671
1090 671
6 0 24 0 0 4096 0 283 0 0 0 4
1240 731
1082 731
1082 706
1086 706
7 0 23 0 0 0 0 283 0 0 0 5
1240 740
1179 740
1179 761
1086 761
1086 745
8 0 22 0 0 12288 0 283 0 0 0 5
1240 749
1198 749
1198 791
1084 791
1084 782
1 5 66 0 0 8320 0 6 79 0 0 4
1823 866
1762 866
1762 651
1804 651
1 6 67 0 0 8320 0 7 79 0 0 4
1823 900
1773 900
1773 660
1804 660
1 7 68 0 0 8320 0 5 79 0 0 4
1823 942
1783 942
1783 669
1804 669
0 0 69 0 0 4224 0 0 0 0 0 4
1877 553
1877 543
1880 543
1880 553
0 0 5 0 0 0 0 0 0 484 484 2
1692 381
1685 381
0 0 13 0 0 0 0 0 0 260 442 4
223 1352
254 1352
254 1276
223 1276
0 0 10 0 0 0 0 0 0 254 249 3
114 386
151 386
151 304
0 0 8 0 0 0 0 0 0 479 171 5
57 338
74 338
74 258
88 258
88 208
0 0 7 0 0 0 0 0 0 255 477 5
28 325
7 325
7 81
84 81
84 108
0 0 61 0 0 4096 0 0 0 472 157 4
537 1521
537 1807
736 1807
736 1887
2 3 2 0 0 0 0 79 79 0 0 4
1798 624
1782 624
1782 633
1798 633
1 0 2 0 0 0 0 79 0 0 211 4
1804 615
1787 615
1787 590
1895 590
10 0 2 0 0 0 0 79 0 0 211 3
1874 624
1895 624
1895 614
12 0 70 0 0 0 0 282 0 0 200 2
1287 548
1287 548
11 0 71 0 0 0 0 282 0 0 199 2
1287 539
1287 539
14 9 72 0 0 8320 0 77 282 0 0 4
1506 786
1360 786
1360 521
1287 521
13 10 73 0 0 12416 0 77 282 0 0 5
1524 786
1524 822
1348 822
1348 530
1287 530
12 0 71 0 0 12416 0 77 0 0 0 5
1542 786
1542 839
1335 839
1335 539
1284 539
11 0 70 0 0 12416 0 77 0 0 0 5
1560 786
1560 829
1324 829
1324 548
1283 548
10 1 2 0 0 0 0 77 76 0 0 3
1497 716
1475 716
1475 749
11 9 32 0 0 8320 0 283 77 0 0 5
1304 722
1388 722
1388 601
1506 601
1506 722
12 7 31 0 0 4224 0 283 77 0 0 5
1304 731
1431 731
1431 641
1524 641
1524 722
14 3 29 0 0 4224 0 283 77 0 0 5
1304 749
1456 749
1456 690
1560 690
1560 722
6 0 74 0 0 4096 0 77 0 0 208 4
1533 722
1533 694
1532 694
1532 679
4 0 75 0 0 4096 0 77 0 0 209 4
1551 722
1551 694
1550 694
1550 679
11 8 76 0 0 12416 0 79 77 0 0 7
1868 651
1934 651
1934 701
1679 701
1679 608
1515 608
1515 722
12 0 74 0 0 12416 0 79 0 0 205 7
1868 660
1903 660
1903 721
1660 721
1660 629
1532 629
1532 683
13 0 75 0 0 12416 0 79 0 0 0 7
1868 669
1916 669
1916 743
1643 743
1643 639
1550 639
1550 684
14 2 77 0 0 12416 0 79 77 0 0 7
1868 678
1890 678
1890 759
1629 759
1629 654
1569 654
1569 722
1 9 2 0 0 0 0 78 79 0 0 3
1895 578
1895 615
1874 615
0 0 22 0 0 0 0 0 0 473 239 2
443 161
484 161
0 0 23 0 0 0 0 0 0 474 240 2
443 154
483 154
0 0 24 0 0 0 0 0 0 475 241 2
442 146
483 146
0 0 25 0 0 0 0 0 0 476 242 2
442 138
482 138
0 3 6 0 0 16384 0 0 297 482 0 7
2112 814
2112 847
1660 847
1660 813
1189 813
1189 888
1217 888
0 0 27 0 0 0 27 0 0 0 487 3
596 65
596 67
737 67
0 0 78 0 0 4096 0 0 0 225 243 2
867 441
867 420
0 0 79 0 0 4096 0 0 0 226 244 2
836 437
836 418
0 0 78 0 0 4096 0 0 0 598 225 2
867 792
867 770
0 0 79 0 0 0 0 0 0 599 226 2
836 793
836 774
0 0 80 0 0 4096 0 0 0 600 227 2
804 793
804 772
0 0 81 0 0 4096 0 0 0 601 228 2
772 790
772 774
0 2 27 0 0 12288 27 0 171 370 0 4
278 1302
357 1302
357 1470
724 1470
0 0 78 0 0 4096 0 0 0 0 0 2
867 778
867 433
0 0 79 0 0 4096 0 0 0 0 0 2
836 779
836 428
0 0 80 0 0 4096 0 0 0 0 245 2
804 780
804 423
0 0 81 0 0 4096 0 0 0 0 0 2
772 780
772 428
0 15 25 0 0 0 0 0 287 0 0 3
697 715
697 684
690 684
0 16 24 0 0 0 0 0 287 0 0 3
702 718
702 693
690 693
0 17 23 0 0 0 0 0 287 0 0 3
707 716
707 702
690 702
0 18 22 0 0 0 0 0 287 0 0 3
725 715
725 711
690 711
0 0 25 0 0 0 0 0 0 234 527 2
790 684
779 684
0 0 25 0 0 0 0 0 0 0 597 2
787 684
924 684
0 0 24 0 0 4096 0 0 0 0 596 2
790 693
954 693
0 0 23 0 0 4096 0 0 0 0 594 2
788 702
984 702
0 0 22 0 0 4096 0 0 0 0 595 2
791 711
1013 711
0 0 27 0 0 0 27 0 0 0 541 2
278 351
278 297
0 0 22 0 0 4096 0 0 0 0 595 2
460 161
1013 161
0 0 23 0 0 4096 0 0 0 0 594 2
461 154
984 154
0 0 24 0 0 4096 0 0 0 0 596 2
463 146
954 146
0 0 25 0 0 4096 0 0 0 0 597 2
465 138
924 138
0 0 78 0 0 0 0 0 0 0 0 2
867 429
867 130
0 0 79 0 0 0 0 0 0 0 0 2
836 424
836 131
0 0 80 0 0 0 0 0 0 0 0 2
804 429
804 132
0 0 81 0 0 0 0 0 0 228 0 2
772 431
772 132
1 0 27 0 0 0 27 277 0 0 0 4
361 200
278 200
278 67
361 67
1 0 11 0 0 0 0 240 0 0 0 3
174 673
168 673
168 739
0 0 10 0 0 0 0 0 0 251 0 4
151 304
112 304
112 303
68 303
2 1 10 0 0 0 0 278 238 0 0 3
578 318
578 304
178 304
0 1 10 0 0 0 0 0 238 0 0 2
148 304
178 304
0 0 18 0 0 8192 0 0 0 0 256 4
1892 499
1873 499
1873 467
1847 467
0 1 11 0 0 16512 0 0 260 248 0 5
168 731
221 731
221 827
169 827
169 2455
0 1 10 0 0 4224 0 0 259 0 0 2
114 365
114 2585
0 1 7 0 0 4224 0 0 256 0 0 2
28 315
28 2768
0 3 18 0 0 4224 0 0 282 0 0 2
1854 467
1281 467
0 1 5 0 0 8320 0 0 249 0 0 3
1894 381
2671 381
2671 2857
0 1 20 0 0 0 0 0 281 10 0 9
2320 361
2320 366
1750 366
1750 361
1722 361
1722 362
1166 362
1166 485
1137 485
0 1 4 0 0 8320 0 0 247 583 0 3
1712 270
2732 270
2732 3024
0 1 13 0 0 4224 0 0 262 0 0 2
223 1347
223 2339
0 1 12 0 0 4224 0 0 261 0 0 4
196 1197
196 2381
226 2381
226 2458
1 0 34 0 0 0 0 8 0 0 0 2
143 755
143 705
0 0 8 0 0 0 0 0 0 0 0 4
45 240
45 239
69 239
69 217
1 1 82 0 0 4224 0 9 287 0 0 2
626 583
626 630
2 1 82 0 0 0 0 287 287 0 0 2
626 639
626 630
3 2 82 0 0 0 0 287 287 0 0 2
626 648
626 639
4 3 82 0 0 0 0 287 287 0 0 2
626 657
626 648
5 4 82 0 0 0 0 287 287 0 0 2
626 666
626 657
6 5 82 0 0 0 0 287 287 0 0 2
626 675
626 666
1 0 22 0 0 0 0 80 0 0 595 2
1013 1350
1013 1350
1 0 23 0 0 0 0 81 0 0 594 2
984 1350
984 1350
1 0 24 0 0 0 0 82 0 0 596 2
954 1350
954 1350
1 0 25 0 0 0 0 83 0 0 597 2
924 1350
924 1350
1 0 78 0 0 0 0 84 0 0 598 2
867 1350
867 1350
1 0 79 0 0 0 0 85 0 0 599 2
836 1350
836 1350
1 0 80 0 0 0 0 86 0 0 600 2
804 1349
804 1349
1 0 81 0 0 0 0 87 0 0 601 2
772 1349
772 1349
1 0 81 0 0 0 0 88 0 0 601 2
772 980
772 980
1 0 80 0 0 0 0 89 0 0 600 2
804 980
804 980
1 0 79 0 0 0 0 90 0 0 599 2
836 980
836 980
1 0 78 0 0 0 0 91 0 0 598 2
867 980
867 980
1 0 25 0 0 0 0 92 0 0 597 2
924 980
924 980
1 0 24 0 0 0 0 93 0 0 596 2
954 980
954 980
1 0 23 0 0 0 0 94 0 0 594 2
984 980
984 980
1 0 22 0 0 0 0 95 0 0 595 2
1013 979
1013 979
1 0 81 0 0 0 0 96 0 0 228 2
772 604
772 604
1 0 80 0 0 0 0 97 0 0 227 2
804 604
804 604
1 0 79 0 0 0 0 98 0 0 226 2
836 603
836 603
0 0 78 0 0 0 0 0 0 0 225 3
880 598
880 603
867 603
1 0 25 0 0 0 0 99 0 0 597 2
924 604
924 604
1 0 24 0 0 0 0 100 0 0 596 2
954 604
954 604
1 0 23 0 0 0 0 101 0 0 594 2
984 604
984 604
1 0 22 0 0 0 0 102 0 0 595 2
1013 604
1013 604
1 0 22 0 0 0 0 103 0 0 536 2
597 277
597 277
1 0 23 0 0 0 0 104 0 0 537 2
597 259
597 259
1 0 24 0 0 0 0 105 0 0 538 2
597 241
597 241
1 0 25 0 0 0 0 106 0 0 539 2
597 223
597 223
1 0 83 0 0 0 0 107 0 0 588 2
473 277
473 277
1 0 84 0 0 0 0 108 0 0 589 2
473 259
473 259
1 0 85 0 0 0 0 109 0 0 590 2
473 241
473 241
1 0 86 0 0 0 0 110 0 0 587 2
473 223
473 223
0 0 23 0 0 0 0 0 0 0 474 3
321 253
321 254
327 254
0 0 24 0 0 0 0 0 0 0 475 2
304 245
318 245
0 0 25 0 0 0 0 0 0 0 476 2
290 236
309 236
1 0 22 0 0 0 0 111 0 0 532 3
736 349
742 349
742 350
1 0 23 0 0 0 0 112 0 0 533 3
714 331
719 331
719 332
1 0 24 0 0 0 0 113 0 0 534 2
687 312
695 312
1 0 25 0 0 0 0 114 0 0 535 3
663 296
672 296
672 297
0 0 87 0 0 4096 0 0 0 0 559 2
617 432
608 432
0 0 88 0 0 4096 0 0 0 0 540 2
599 423
590 423
0 0 89 0 0 8192 0 0 0 0 561 3
581 413
581 414
571 414
0 0 90 0 0 4096 0 0 0 0 562 2
563 406
548 406
1 0 87 0 0 0 0 115 0 0 559 2
608 621
608 621
1 0 88 0 0 0 0 116 0 0 560 2
590 621
590 621
1 0 89 0 0 0 0 117 0 0 561 2
572 621
572 622
1 0 90 0 0 0 0 118 0 0 562 2
554 621
554 621
1 0 22 0 0 0 0 119 0 0 524 2
759 711
759 711
1 0 23 0 0 0 0 120 0 0 525 2
759 702
759 702
1 0 24 0 0 0 0 121 0 0 526 2
759 693
759 693
1 0 25 0 0 0 0 122 0 0 527 2
759 684
759 684
1 0 78 0 0 0 0 123 0 0 528 2
759 675
759 675
1 0 79 0 0 0 0 124 0 0 529 2
759 666
759 666
1 0 80 0 0 0 0 125 0 0 530 2
759 657
759 657
1 0 81 0 0 0 0 126 0 0 531 2
759 648
759 648
1 0 22 0 0 0 0 127 0 0 516 2
719 1161
719 1161
1 0 23 0 0 0 0 128 0 0 517 2
698 1152
698 1152
1 0 24 0 0 0 0 129 0 0 518 2
679 1143
679 1143
1 0 25 0 0 0 0 130 0 0 519 2
660 1134
660 1134
1 0 78 0 0 0 0 131 0 0 520 2
485 1277
485 1277
1 0 79 0 0 0 0 132 0 0 521 2
471 1267
471 1267
1 0 80 0 0 0 0 133 0 0 522 2
460 1258
460 1258
1 0 81 0 0 0 0 134 0 0 523 2
449 1248
449 1248
1 0 60 0 0 0 0 135 0 0 469 2
510 1343
510 1343
1 0 63 0 0 0 0 136 0 0 470 2
519 1322
519 1322
1 0 62 0 0 0 0 137 0 0 471 2
528 1301
528 1301
1 0 61 0 0 0 0 138 0 0 472 2
538 1285
537 1285
1 0 22 0 0 0 0 139 0 0 546 2
742 1113
742 1113
1 0 23 0 0 0 0 140 0 0 547 2
735 1104
735 1104
1 0 24 0 0 0 0 141 0 0 548 2
724 1095
724 1095
1 0 25 0 0 0 0 142 0 0 549 2
711 1086
711 1086
1 0 22 0 0 0 0 143 0 0 512 2
1060 345
1060 345
1 0 23 0 0 0 0 144 0 0 513 2
1060 327
1060 327
1 0 24 0 0 0 0 145 0 0 514 2
1060 309
1060 309
1 0 25 0 0 0 0 146 0 0 515 2
1060 291
1060 291
1 0 17 0 0 0 0 147 0 0 579 2
1184 346
1184 345
1 0 14 0 0 0 0 148 0 0 580 2
1184 327
1184 327
1 0 16 0 0 0 0 149 0 0 581 2
1184 309
1184 309
1 0 15 0 0 0 0 150 0 0 582 2
1183 291
1183 291
1 0 91 0 0 0 0 151 0 0 572 2
1160 548
1160 548
1 0 92 0 0 0 0 152 0 0 573 2
1160 530
1160 530
1 0 93 0 0 0 0 153 0 0 574 2
1160 512
1160 512
1 0 94 0 0 0 0 154 0 0 575 2
1160 494
1160 494
1 0 17 0 0 0 0 155 0 0 568 2
1349 413
1349 413
1 0 14 0 0 0 0 156 0 0 569 2
1335 413
1335 413
1 0 16 0 0 0 0 157 0 0 570 2
1321 413
1321 413
1 0 15 0 0 0 0 158 0 0 571 2
1308 413
1308 413
1 0 17 0 0 0 0 159 0 0 579 2
1349 231
1349 231
1 0 14 0 0 0 0 160 0 0 580 2
1335 231
1335 231
1 0 16 0 0 0 0 161 0 0 581 2
1321 231
1321 231
1 0 15 0 0 0 0 162 0 0 582 2
1308 231
1308 231
1 0 22 0 0 0 0 163 0 0 492 2
1114 933
1114 933
1 0 23 0 0 0 0 164 0 0 493 2
1093 924
1093 924
1 0 24 0 0 0 0 165 0 0 494 2
1070 915
1070 915
1 0 25 0 0 0 0 166 0 0 495 2
1050 905
1050 906
1 0 22 0 0 0 0 167 0 0 504 2
1110 224
1110 224
1 0 23 0 0 0 0 168 0 0 505 2
1086 215
1086 215
1 0 24 0 0 0 0 169 0 0 506 2
1061 206
1061 206
1 0 25 0 0 0 0 170 0 0 507 2
1040 197
1040 197
1 3 95 0 0 4224 0 171 273 0 0 2
758 1470
1176 1470
4 0 27 0 0 8320 27 288 0 0 0 4
439 1191
278 1191
278 2307
327 2307
1 0 3 0 0 0 0 172 0 0 481 2
2761 3083
2761 3083
1 0 4 0 0 0 0 173 0 0 259 2
2732 2996
2732 2996
1 0 5 0 0 0 0 175 0 0 257 2
2671 2838
2671 2838
1 0 5 0 0 0 0 180 0 0 483 2
2522 2466
2522 2466
1 0 6 0 0 0 0 181 0 0 482 2
2463 2308
2464 2308
1 0 3 0 0 0 0 182 0 0 481 2
2762 2276
2761 2276
1 0 4 0 0 0 0 183 0 0 259 2
2731 2254
2732 2254
1 0 5 0 0 0 0 185 0 0 257 2
2671 2206
2671 2206
1 0 5 0 0 0 0 186 0 0 483 2
2522 2092
2522 2092
1 0 6 0 0 0 0 187 0 0 482 2
2463 2036
2464 2036
1 0 3 0 0 0 0 188 0 0 481 2
2761 1748
2761 1748
1 0 4 0 0 0 0 189 0 0 259 2
2732 1732
2732 1732
1 0 5 0 0 0 0 190 0 0 257 2
2670 1696
2671 1696
1 0 5 0 0 0 0 191 0 0 483 2
2522 1616
2522 1616
1 0 6 0 0 0 0 192 0 0 386 2
2463 1549
2463 1549
1 0 6 0 0 0 0 193 0 0 482 2
2463 1549
2464 1549
1 0 3 0 0 0 0 194 0 0 481 2
2762 1325
2761 1325
1 0 4 0 0 0 0 195 0 0 259 2
2733 1304
2732 1304
1 0 5 0 0 0 0 196 0 0 257 2
2671 1269
2671 1269
1 0 5 0 0 0 0 197 0 0 483 2
2522 1170
2522 1170
1 0 6 0 0 0 0 198 0 0 482 2
2463 1131
2464 1131
1 0 3 0 0 0 0 199 0 0 481 2
2761 562
2761 562
1 0 4 0 0 0 0 200 0 0 259 2
2732 538
2732 538
1 0 5 0 0 0 0 201 0 0 257 2
2671 488
2671 488
1 0 5 0 0 0 0 202 0 0 483 2
2522 523
2522 523
1 0 3 0 0 0 0 203 0 0 481 2
2761 921
2761 921
1 0 4 0 0 0 0 204 0 0 259 2
2732 900
2732 900
1 0 5 0 0 0 0 205 0 0 257 2
2671 865
2671 865
1 0 5 0 0 0 0 206 0 0 483 2
2522 750
2522 750
1 0 7 0 0 0 0 207 0 0 255 2
27 2756
28 2756
1 0 8 0 0 0 0 208 0 0 479 2
57 2698
57 2698
1 0 9 0 0 0 0 209 0 0 480 2
85 2634
86 2634
1 0 10 0 0 0 0 210 0 0 254 2
113 2570
114 2570
1 0 11 0 0 0 0 211 0 0 253 2
169 2442
169 2442
1 0 12 0 0 0 0 212 0 0 261 2
196 2381
196 2381
1 0 13 0 0 0 0 213 0 0 260 2
223 2327
223 2327
1 0 13 0 0 0 0 214 0 0 260 2
224 2062
223 2062
1 0 12 0 0 0 0 215 0 0 261 2
196 2015
196 2015
1 0 11 0 0 0 0 216 0 0 253 2
169 1967
169 1967
1 0 10 0 0 0 0 217 0 0 254 2
113 1850
114 1850
1 0 9 0 0 0 0 218 0 0 480 2
86 1794
86 1794
1 0 8 0 0 0 0 219 0 0 479 2
57 1744
57 1744
1 0 7 0 0 0 0 220 0 0 255 2
28 1704
28 1704
1 0 13 0 0 0 0 221 0 0 260 2
223 1450
223 1450
1 0 12 0 0 0 0 222 0 0 261 2
196 1394
196 1394
1 0 11 0 0 0 0 223 0 0 253 2
169 1348
169 1348
1 0 10 0 0 0 0 224 0 0 254 2
115 1266
114 1266
1 0 9 0 0 0 0 225 0 0 480 2
85 1230
86 1230
1 0 8 0 0 0 0 226 0 0 479 2
57 1184
57 1184
1 0 7 0 0 0 0 227 0 0 255 2
28 1140
28 1140
1 0 13 0 0 0 0 228 0 0 442 2
223 1191
223 1191
1 0 12 0 0 0 0 229 0 0 441 2
196 1026
196 1026
1 0 11 0 0 0 0 230 0 0 253 2
169 924
169 924
1 0 10 0 0 0 0 231 0 0 254 2
114 842
114 842
1 0 9 0 0 0 0 232 0 0 480 2
86 788
86 788
1 0 8 0 0 0 0 233 0 0 479 2
57 749
57 749
1 0 7 0 0 0 0 234 0 0 255 2
28 725
28 725
0 0 10 0 0 0 0 0 0 0 254 3
149 531
149 536
114 536
0 0 8 0 0 0 0 0 0 0 479 2
69 448
57 448
0 0 7 0 0 0 0 0 0 0 255 3
40 415
40 414
28 414
1 0 7 0 0 0 0 235 0 0 477 4
517 108
516 108
516 109
515 109
1 0 7 0 0 0 0 236 0 0 477 2
179 107
179 108
1 0 8 0 0 0 0 237 0 0 171 2
144 209
144 208
1 0 34 0 0 0 0 239 0 0 161 2
174 644
174 644
0 0 6 0 0 0 0 0 0 0 216 3
1648 862
1648 813
1634 813
1 0 18 0 0 0 0 242 0 0 256 2
1707 467
1707 467
1 0 2 0 0 0 0 244 0 0 168 2
1625 448
1625 449
0 0 96 0 0 4096 0 0 0 0 485 3
1634 414
1634 401
1625 401
0 0 20 0 0 0 0 0 0 0 258 3
1622 343
1622 362
1625 362
1 0 4 0 0 0 0 245 0 0 583 2
1622 269
1622 270
9 0 12 0 0 0 0 291 0 0 172 5
713 1050
714 1050
714 1026
196 1026
196 1092
2 0 13 0 0 0 0 288 0 0 0 3
433 1173
223 1173
223 1282
1 0 7 0 0 0 0 263 0 0 464 2
911 1627
911 1627
1 0 8 0 0 0 0 264 0 0 463 2
911 1654
911 1654
1 0 40 0 0 0 0 265 0 0 448 2
911 1684
911 1684
1 0 58 0 0 0 0 266 0 0 462 2
911 1712
911 1712
0 1 97 0 0 4096 0 0 11 459 0 2
1168 1528
1069 1528
9 1 40 0 0 20608 0 273 268 0 0 6
1246 1461
1263 1461
1263 1599
798 1599
798 1684
2272 1684
12 2 98 0 0 12416 0 272 273 0 0 6
1477 1503
1521 1503
1521 1240
1118 1240
1118 1461
1182 1461
11 1 8 0 0 0 0 272 273 0 0 6
1471 1494
1512 1494
1512 1272
1128 1272
1128 1452
1182 1452
10 5 7 0 0 0 0 272 272 0 0 6
1477 1467
1484 1467
1484 1409
1373 1409
1373 1485
1407 1485
9 6 99 0 0 16512 0 272 272 0 0 6
1471 1458
1493 1458
1493 1309
1364 1309
1364 1494
1407 1494
12 1 100 0 0 12416 0 273 272 0 0 4
1252 1506
1327 1506
1327 1449
1407 1449
11 2 58 0 0 0 0 273 272 0 0 4
1246 1497
1335 1497
1335 1458
1407 1458
10 6 101 0 0 16512 0 273 273 0 0 6
1252 1470
1271 1470
1271 1318
1146 1318
1146 1497
1182 1497
9 5 40 0 0 0 0 273 273 0 0 6
1246 1461
1263 1461
1263 1352
1155 1352
1155 1488
1182 1488
3 0 95 0 0 0 0 273 0 0 466 5
1176 1470
1175 1470
1175 1432
1398 1432
1398 1468
7 3 95 0 0 0 0 273 273 0 0 4
1176 1506
1175 1506
1175 1470
1176 1470
8 8 97 0 0 12416 0 273 272 0 0 6
1176 1515
1168 1515
1168 1528
1390 1528
1390 1512
1401 1512
8 4 97 0 0 0 0 272 272 0 0 4
1401 1512
1390 1512
1390 1476
1401 1476
4 8 97 0 0 0 0 273 273 0 0 4
1176 1479
1168 1479
1168 1515
1176 1515
11 1 58 0 0 20608 0 273 267 0 0 6
1246 1497
1291 1497
1291 1608
809 1608
809 1712
2273 1712
11 1 8 0 0 20480 0 272 269 0 0 6
1471 1494
1512 1494
1512 1588
786 1588
786 1654
2272 1654
10 1 7 0 0 0 0 272 270 0 0 6
1477 1467
1484 1467
1484 1579
776 1579
776 1627
2272 1627
1 0 95 0 0 0 0 271 0 0 369 2
1025 1452
1025 1470
7 3 95 0 0 0 0 272 272 0 0 4
1401 1503
1398 1503
1398 1467
1401 1467
1 0 27 0 0 0 27 274 0 0 468 2
221 50
221 67
0 3 27 0 0 0 27 0 275 247 0 4
279 67
221 67
221 64
182 64
14 0 60 0 0 8320 0 288 0 0 160 5
503 1227
510 1227
510 1759
763 1759
763 1860
13 0 63 0 0 8320 0 288 0 0 159 5
503 1218
519 1218
519 1775
754 1775
754 1869
12 0 62 0 0 8320 0 288 0 0 0 3
503 1209
528 1209
528 1666
11 0 61 0 0 8320 0 288 0 0 0 3
503 1200
537 1200
537 1528
8 0 22 0 0 0 0 277 0 0 0 4
361 263
335 263
335 161
456 161
7 0 23 0 0 0 0 277 0 0 0 4
361 254
327 254
327 154
457 154
6 0 24 0 0 0 0 277 0 0 0 4
361 245
318 245
318 146
459 146
5 0 25 0 0 0 0 277 0 0 0 4
361 236
309 236
309 138
461 138
1 0 7 0 0 0 0 276 0 0 0 5
526 214
515 214
515 108
50 108
50 109
4 1 102 0 0 4224 0 277 10 0 0 4
361 227
261 227
261 262
260 262
1 0 8 0 0 4224 0 257 0 0 0 2
57 2705
57 319
1 0 9 0 0 4224 0 258 0 0 0 2
86 2647
86 732
1 0 3 0 0 4224 0 246 0 0 0 3
2761 3106
2761 108
1853 108
1 0 6 0 0 4224 0 255 0 0 0 3
2464 2322
2464 814
2098 814
1 0 5 0 0 0 0 254 0 0 0 3
2522 2482
2522 476
2056 476
14 0 5 0 0 0 0 282 0 0 0 5
1217 458
1204 458
1204 381
1716 381
1716 382
13 1 96 0 0 12416 0 282 1 0 0 6
1217 449
1213 449
1213 401
1716 401
1716 401
1715 401
0 0 27 0 0 0 27 0 0 554 238 2
278 1077
278 321
0 0 27 0 0 0 27 0 0 489 0 2
1146 67
725 67
0 4 27 0 0 0 27 0 297 489 0 5
1417 564
1417 797
1176 797
1176 897
1223 897
4 4 27 0 0 0 27 279 283 0 0 8
1221 188
1146 188
1146 67
1417 67
1417 564
1175 564
1175 713
1240 713
0 0 24 0 0 0 0 0 0 596 0 2
954 512
1014 512
0 0 25 0 0 0 0 0 0 597 19 2
924 494
1064 494
8 0 22 0 0 0 0 297 0 0 595 2
1223 933
1013 933
7 0 23 0 0 0 0 297 0 0 594 2
1223 924
984 924
6 0 24 0 0 0 0 297 0 0 596 2
1223 915
954 915
5 0 25 0 0 0 0 297 0 0 597 2
1223 906
924 906
14 1 103 0 0 4224 0 297 293 0 0 4
1287 933
1444 933
1444 896
1443 896
13 1 104 0 0 4224 0 297 292 0 0 3
1287 924
1420 924
1420 896
12 1 105 0 0 4224 0 297 294 0 0 3
1287 915
1397 915
1397 896
11 1 106 0 0 4224 0 297 295 0 0 3
1287 906
1374 906
1374 896
9 1 2 0 0 0 0 297 296 0 0 2
1293 870
1293 846
3 2 6 0 0 0 0 297 297 0 0 2
1217 888
1217 879
10 9 2 0 0 0 0 297 297 0 0 2
1293 879
1293 870
1 9 2 0 0 0 0 297 297 0 0 5
1223 870
1213 870
1213 850
1293 850
1293 870
8 0 22 0 0 0 0 279 0 0 595 2
1221 224
1013 224
7 0 23 0 0 0 0 279 0 0 594 2
1221 215
984 215
6 0 24 0 0 0 0 279 0 0 596 2
1221 206
954 206
5 0 25 0 0 0 0 279 0 0 597 2
1221 197
924 197
10 1 2 0 0 0 0 279 285 0 0 4
1291 170
1301 170
1301 170
1298 170
3 2 3 0 0 0 0 279 279 0 0 2
1215 179
1215 170
10 9 2 0 0 0 0 279 279 0 0 2
1291 170
1291 161
1 9 2 0 0 0 0 279 279 0 0 5
1221 161
1220 161
1220 141
1291 141
1291 161
12 0 22 0 0 0 0 280 0 0 595 2
1071 345
1013 345
11 0 23 0 0 0 0 280 0 0 594 2
1071 327
984 327
10 0 24 0 0 0 0 280 0 0 596 2
1071 309
954 309
9 0 25 0 0 0 0 280 0 0 597 2
1071 291
924 291
8 0 22 0 0 0 0 291 0 0 595 4
643 1113
618 1113
618 1161
1013 1161
7 0 23 0 0 0 0 291 0 0 594 4
643 1104
609 1104
609 1152
984 1152
6 0 24 0 0 0 0 291 0 0 596 4
643 1095
600 1095
600 1143
954 1143
5 0 25 0 0 0 0 291 0 0 597 4
643 1086
591 1086
591 1134
924 1134
8 0 78 0 0 12288 0 288 0 0 598 4
439 1227
418 1227
418 1277
867 1277
7 0 79 0 0 12288 0 288 0 0 599 4
439 1218
407 1218
407 1267
836 1267
6 0 80 0 0 12288 0 288 0 0 600 4
439 1209
397 1209
397 1258
804 1258
5 0 81 0 0 12288 0 288 0 0 601 4
439 1200
387 1200
387 1248
772 1248
18 0 22 0 0 0 0 287 0 0 237 2
690 711
794 711
17 0 23 0 0 0 0 287 0 0 236 2
690 702
792 702
16 0 24 0 0 0 0 287 0 0 235 2
690 693
793 693
15 0 25 0 0 0 0 287 0 0 0 2
690 684
783 684
14 0 78 0 0 0 0 287 0 0 225 2
690 675
867 675
13 0 79 0 0 0 0 287 0 0 226 2
690 666
836 666
12 0 80 0 0 0 0 287 0 0 227 2
690 657
804 657
11 0 81 0 0 0 0 287 0 0 228 2
690 648
772 648
8 0 22 0 0 0 0 278 0 0 595 4
632 324
650 324
650 350
1013 350
7 0 23 0 0 0 0 278 0 0 594 5
623 324
623 319
657 319
657 332
984 332
6 0 24 0 0 0 0 278 0 0 596 3
614 324
614 312
954 312
5 0 25 0 0 0 0 278 0 0 597 3
605 324
605 297
924 297
12 0 22 0 0 0 0 276 0 0 595 2
590 277
1013 277
11 0 23 0 0 0 0 276 0 0 594 2
590 259
984 259
10 0 24 0 0 0 0 276 0 0 596 2
590 241
954 241
9 0 25 0 0 0 0 276 0 0 597 2
590 223
924 223
0 13 88 0 0 4096 0 0 278 560 0 4
590 560
590 423
623 423
623 388
4 0 27 0 0 0 27 278 0 0 0 4
596 324
596 297
278 297
278 261
2 3 10 0 0 0 0 278 278 0 0 2
578 318
587 318
1 1 2 0 0 0 0 278 284 0 0 3
569 324
569 323
541 323
1 9 2 0 0 0 0 278 278 0 0 5
569 324
569 323
546 323
546 394
569 394
10 9 2 0 0 0 0 278 278 0 0 2
578 394
569 394
14 0 22 0 0 0 0 291 0 0 595 2
707 1113
1013 1113
13 0 23 0 0 0 0 291 0 0 594 2
707 1104
984 1104
12 0 24 0 0 0 0 291 0 0 596 2
707 1095
954 1095
11 0 25 0 0 0 0 291 0 0 597 2
707 1086
924 1086
1 1 2 0 0 0 0 291 290 0 0 3
643 1050
627 1050
627 1044
3 2 13 0 0 0 0 291 288 0 0 5
637 1068
637 1059
422 1059
422 1173
433 1173
3 2 13 0 0 0 0 291 291 0 0 2
637 1068
637 1059
10 9 12 0 0 0 0 291 291 0 0 4
713 1059
714 1059
714 1050
713 1050
4 4 27 0 0 0 27 291 288 0 0 4
643 1077
278 1077
278 1191
439 1191
9 1 2 0 0 0 0 288 289 0 0 4
509 1164
524 1164
524 1164
519 1164
3 2 13 0 0 0 0 288 288 0 0 4
433 1182
422 1182
422 1173
433 1173
10 9 2 0 0 0 0 288 288 0 0 4
509 1173
510 1173
510 1164
509 1164
1 9 2 0 0 0 0 288 288 0 0 6
439 1164
438 1164
438 1144
510 1144
510 1164
509 1164
10 14 87 0 0 8320 0 287 278 0 0 5
626 711
608 711
608 432
632 432
632 388
9 0 88 0 0 8320 0 287 0 0 540 3
626 702
590 702
590 554
8 12 89 0 0 8320 0 287 278 0 0 7
626 693
572 693
572 519
571 519
571 414
614 414
614 388
7 11 90 0 0 8320 0 287 278 0 0 7
626 684
554 684
554 529
548 529
548 405
605 405
605 388
19 1 11 0 0 0 0 287 240 0 0 6
696 630
700 630
700 600
511 600
511 673
174 673
9 1 2 0 0 0 0 283 286 0 0 5
1310 686
1291 686
1291 617
1284 617
1284 613
3 2 33 0 0 0 0 283 283 0 0 7
1234 704
1224 704
1224 650
1216 650
1216 650
1234 650
1234 695
10 9 2 0 0 0 0 283 283 0 0 4
1310 695
1310 641
1310 641
1310 686
1 9 2 0 0 0 0 283 283 0 0 5
1240 686
1212 686
1212 617
1310 617
1310 686
0 8 17 0 0 0 0 0 282 579 0 3
1349 345
1349 512
1287 512
0 7 14 0 0 0 0 0 282 580 0 3
1335 327
1335 503
1287 503
0 6 16 0 0 0 0 0 282 581 0 3
1321 309
1321 494
1287 494
0 5 15 0 0 0 0 0 282 582 0 3
1308 291
1308 485
1287 485
8 22 91 0 0 4224 0 281 282 0 0 2
1137 548
1211 548
6 21 92 0 0 4224 0 281 282 0 0 4
1137 530
1184 530
1184 539
1211 539
20 4 93 0 0 12416 0 282 281 0 0 4
1211 530
1195 530
1195 512
1137 512
2 19 94 0 0 4224 0 281 282 0 0 4
1137 494
1206 494
1206 521
1211 521
5 7 20 0 0 0 0 281 281 0 0 4
1137 521
1166 521
1166 539
1137 539
3 5 20 0 0 0 0 281 281 0 0 4
1137 503
1166 503
1166 521
1137 521
1 3 20 0 0 0 0 281 281 0 0 4
1137 485
1166 485
1166 503
1137 503
8 14 17 0 0 0 0 280 279 0 0 4
1135 345
1349 345
1349 224
1285 224
6 13 14 0 0 0 0 280 279 0 0 4
1135 327
1335 327
1335 215
1285 215
4 12 16 0 0 0 0 280 279 0 0 4
1135 309
1321 309
1321 206
1285 206
2 11 15 0 0 0 0 280 279 0 0 4
1135 291
1308 291
1308 197
1285 197
1 0 4 0 0 0 0 280 0 0 0 4
1135 282
1144 282
1144 270
1725 270
5 7 4 0 0 0 0 280 280 0 0 4
1135 318
1144 318
1144 336
1135 336
3 5 4 0 0 0 0 280 280 0 0 4
1135 300
1144 300
1144 318
1135 318
1 3 4 0 0 0 0 280 280 0 0 4
1135 282
1144 282
1144 300
1135 300
11 2 86 0 0 12416 0 277 276 0 0 4
425 236
458 236
458 223
526 223
14 8 83 0 0 12416 0 277 276 0 0 4
425 263
457 263
457 277
526 277
13 6 84 0 0 12416 0 277 276 0 0 4
425 254
468 254
468 259
526 259
12 4 85 0 0 12416 0 277 276 0 0 4
425 245
468 245
468 241
526 241
7 5 7 0 0 0 0 276 276 0 0 4
526 268
515 268
515 250
526 250
5 3 7 0 0 0 0 276 276 0 0 4
526 250
515 250
515 232
526 232
3 1 7 0 0 0 0 276 276 0 0 4
526 232
515 232
515 214
526 214
0 0 23 0 0 4224 0 0 0 0 0 2
984 1369
984 128
0 1 22 0 0 4224 0 0 0 0 0 2
1013 1369
1013 126
0 0 24 0 0 4224 0 0 0 0 0 2
954 1369
954 129
0 0 25 0 0 4224 0 0 0 0 0 2
924 1369
924 130
0 0 78 0 0 4224 0 0 0 0 0 2
867 1369
867 782
0 0 79 0 0 4224 0 0 0 0 0 2
836 1369
836 783
0 0 80 0 0 4224 0 0 0 0 0 2
804 1369
804 784
0 0 81 0 0 4224 0 0 0 0 0 2
772 1369
772 784
148
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1086 1802 1111 1846
1094 1810 1102 1842
5 T
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1153 2118 1222 2142
1163 2126 1211 2142
6 lda t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
1464 2349 1492 2416
1474 2359 1481 2414
18 C
e 
b
a
r
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2480 2636 2523 2651
2494 2647 2508 2658
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2414 2599 2459 2614
2429 2610 2443 2621
2 Zf
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
2316 2527 2394 2542
2330 2539 2379 2550
7 Se S3 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1882 2429 1949 2444
1897 2440 1933 2451
5 Jz t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2176 2601 2219 2616
2190 2613 2204 2624
2 Lo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2066 2636 2109 2651
2080 2647 2094 2658
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1940 2630 2010 2645
1954 2641 1995 2652
6 lb bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1800 2631 1870 2646
1814 2643 1855 2654
6 Ei bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1669 2610 1739 2625
1683 2621 1724 2632
6 la bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1761 2369 1828 2384
1776 2380 1812 2391
5 xr t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1649 2367 1719 2382
1663 2379 1704 2390
6 sub t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1319 2259 1389 2274
1333 2270 1374 2281
6 Li bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1229 2270 1272 2285
1243 2281 1257 2292
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1150 2298 1219 2322
1160 2306 1208 2322
6 lm bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1060 2133 1097 2157
1070 2141 1086 2157
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
359 1896 476 1920
369 1904 465 1920
12 control unit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1116 654 1149 678
1124 662 1140 678
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1118 770 1151 794
1126 778 1142 794
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1849 849 1882 873
1857 857 1873 873
2 C3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1837 986 1870 1010
1845 994 1861 1010
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1215 586 1276 610
1225 594 1265 610
5 B REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1807 563 1868 587
1817 571 1857 587
5 C REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
911 105 944 129
919 113 935 129
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
415 281 454 305
422 286 446 302
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
201 210 264 234
208 216 256 232
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
278 1444 317 1468
285 1449 309 1465
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
701 592 764 616
708 598 756 614
6 WE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1162 105 1225 129
1169 110 1217 126
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
472 1405 575 1429
479 1411 567 1427
11 I4 I5 I6 I7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1288 1541 1319 1565
1295 1547 1311 1563
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1239 1541 1270 1565
1246 1547 1262 1563
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1508 1531 1539 1555
1515 1536 1531 1552
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1164 247 1195 271
1171 253 1187 269
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1140 366 1171 390
1147 371 1163 387
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
482 84 513 108
489 89 505 105
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
226 85 257 109
233 90 249 106
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
216 190 247 214
223 195 239 211
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
273 875 312 899
280 880 304 896
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1454 788 1517 812
1461 793 1509 809
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 462 1478 486
1454 468 1470 484
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 452 1478 476
1454 458 1470 474
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 442 1478 466
1454 448 1470 464
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 433 1478 457
1454 439 1470 455
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1452 382 1491 406
1459 388 1483 404
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1490 362 1513 386
1497 368 1505 384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
213 1143 276 1167
220 1149 268 1165
6 Li BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
217 996 280 1020
224 1001 272 1017
6 Ei BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
208 647 271 671
215 653 263 669
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
208 617 271 641
215 623 263 639
6 WE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
200 280 263 304
207 286 255 302
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
277 1168 316 1192
284 1173 308 1189
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
272 1053 311 1077
279 1058 303 1074
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
878 43 917 67
885 48 909 64
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
275 64 314 88
282 69 306 85
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1376 769 1415 793
1383 774 1407 790
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1378 539 1417 563
1385 544 1409 560
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1367 44 1406 68
1374 49 1398 65
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
639 563 678 587
646 569 670 585
3 RAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
852 108 883 132
859 113 875 129
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
820 109 851 133
827 114 843 130
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 109 819 133
795 114 811 130
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
757 108 788 132
764 114 780 130
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
999 107 1030 131
1006 113 1022 129
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
969 107 1000 131
976 113 992 129
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
938 108 969 132
945 113 961 129
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1232 410 1275 431
1241 416 1265 431
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1235 114 1270 138
1240 118 1264 134
3 ACC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
650 361 685 385
655 365 679 381
3 MAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
380 161 407 185
385 165 401 181
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1214 817 1285 841
1221 822 1277 838
7 O/P REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
818 1608 849 1632
825 1613 841 1629
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
817 1634 848 1658
824 1639 840 1655
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
818 1661 849 1685
825 1667 841 1683
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
818 1690 849 1714
825 1696 841 1712
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2306 1699 2337 1723
2313 1705 2329 1721
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2306 1672 2337 1696
2313 1678 2329 1694
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2305 1646 2336 1670
2312 1651 2328 1667
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2303 1616 2334 1640
2310 1621 2326 1637
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2378 787 2441 811
2385 792 2433 808
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 473 2537 497
2513 479 2529 495
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1787 453 1818 477
1794 459 1810 475
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1816 462 1847 486
1823 468 1839 484
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1763 444 1794 468
1770 450 1786 466
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1736 435 1767 459
1743 441 1759 457
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2178 462 2209 486
2185 468 2201 484
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1911 382 1950 406
1918 388 1942 404
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1953 362 1976 386
1960 368 1968 384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2332 362 2355 386
2339 368 2347 384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2293 382 2332 406
2300 388 2324 404
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 436 2683 460
2667 442 2675 458
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1190 377 1213 401
1197 383 1205 399
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1208 394 1247 418
1215 400 1239 416
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2368 250 2399 274
2375 256 2391 272
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2708 249 2739 273
2715 255 2731 271
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2371 88 2434 112
2378 93 2426 109
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2705 89 2768 113
2712 94 2760 110
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2507 743 2538 767
2514 749 2530 765
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1017 2537 1041
2513 1023 2529 1039
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1284 2537 1308
2513 1290 2529 1306
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1612 2537 1636
2513 1618 2529 1634
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1932 2537 1956
2513 1938 2529 1954
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2507 2219 2538 2243
2514 2225 2530 2241
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 486 2748 510
2724 492 2740 508
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2737 290 2800 314
2744 295 2792 311
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2736 510 2799 534
2743 515 2791 531
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 859 2683 883
2667 865 2675 881
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 1098 2683 1122
2667 1104 2675 1120
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 1362 2683 1386
2667 1368 2675 1384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 893 2748 917
2724 899 2740 915
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2736 913 2799 937
2743 918 2791 934
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 1392 2748 1416
2724 1398 2740 1414
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 1693 2683 1717
2667 1699 2675 1715
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 1723 2748 1747
2724 1729 2740 1745
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2738 1743 2801 1767
2745 1748 2793 1764
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 2022 2683 2046
2667 2028 2675 2044
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 2312 2683 2336
2667 2318 2675 2334
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2689 2041 2720 2065
2696 2046 2712 2062
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2689 2331 2720 2355
2696 2336 2712 2352
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 2061 2748 2085
2724 2067 2740 2083
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 2351 2748 2375
2724 2357 2740 2373
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2738 2081 2801 2105
2745 2086 2793 2102
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2737 2374 2800 2398
2744 2379 2792 2395
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2736 2795 2799 2819
2743 2800 2791 2816
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2716 2723 2747 2747
2723 2729 2739 2745
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 2597 2683 2621
2667 2603 2675 2619
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2624 2511 2663 2535
2631 2517 2655 2533
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2596 2462 2627 2486
2603 2468 2619 2484
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 2425 2599 2446
2574 2432 2590 2447
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2433 947 2496 971
2440 952 2488 968
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2433 1215 2496 1239
2440 1220 2488 1236
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2434 1548 2497 1572
2441 1553 2489 1569
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2435 1877 2498 1901
2442 1882 2490 1898
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2434 2153 2497 2177
2441 2158 2489 2174
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
143 2189 206 2213
150 2195 198 2211
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
89 2286 152 2310
96 2292 144 2308
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
61 2348 124 2372
68 2354 116 2370
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 2402 75 2426
51 2407 67 2423
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 2460 45 2484
21 2465 37 2481
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1572 781 1617 805
1582 789 1606 805
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1515 545 1584 569
1525 553 1573 569
6 Lc BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
2271 1737 2380 1761
2281 1745 2369 1761
11 LDAM (0000)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2826 766 2896 781
2840 777 2881 788
6 lb Bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1450 493 1520 508
1464 504 1505 515
6 lb Bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1036 1536 1137 1580
1047 1544 1125 1576
13 must be hight
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
442 1089 489 1153
453 1098 477 1146
10   IR
 MSB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
