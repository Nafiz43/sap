CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
28 D:\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
390
13 Logic Switch~
5 690 1510 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V37
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3713 0 0
2
43746 0
0
13 Logic Switch~
5 457 1892 0 1 11
0 48
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V35
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4635 0 0
2
5.89911e-315 0
0
13 Logic Switch~
5 481 1881 0 1 11
0 49
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V34
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4444 0 0
2
5.89911e-315 5.26354e-315
0
13 Logic Switch~
5 501 1871 0 1 11
0 50
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V24
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3328 0 0
2
5.89911e-315 5.30499e-315
0
13 Logic Switch~
5 527 1860 0 1 11
0 47
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V23
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
312 0 0
2
5.89911e-315 5.32571e-315
0
13 Logic Switch~
5 499 56 0 1 11
0 53
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V32
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8412 0 0
2
43746 1
0
13 Logic Switch~
5 472 735 0 1 11
0 54
0
0 0 20848 90
2 0V
11 -5 25 3
3 V28
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6185 0 0
2
43746 2
0
13 Logic Switch~
5 1817 1001 0 1 11
0 62
0
0 0 20848 180
2 0V
-7 -16 7 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6455 0 0
2
5.89911e-315 5.34643e-315
0
13 Logic Switch~
5 1104 671 0 1 11
0 63
0
0 0 20848 180
2 0V
-7 -16 7 -8
3 V46
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3265 0 0
2
5.89911e-315 5.3568e-315
0
13 Logic Switch~
5 1100 706 0 1 11
0 64
0
0 0 20848 180
2 0V
-7 -16 7 -8
3 V45
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9479 0 0
2
5.89911e-315 5.36716e-315
0
13 Logic Switch~
5 1100 745 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 20848 180
2 5V
-7 -16 7 -8
3 V44
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9330 0 0
2
5.89911e-315 5.37752e-315
0
13 Logic Switch~
5 1098 782 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 20848 180
2 5V
-7 -16 7 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6531 0 0
2
5.89911e-315 5.38788e-315
0
13 Logic Switch~
5 1837 942 0 1 11
0 69
0
0 0 20848 180
2 0V
-7 -16 7 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9789 0 0
2
5.89911e-315 5.39306e-315
0
13 Logic Switch~
5 1837 866 0 10 11
0 67 0 0 0 0 0 0 0 0
1
0
0 0 20848 180
2 5V
-7 -16 7 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8535 0 0
2
5.89911e-315 5.39824e-315
0
13 Logic Switch~
5 1837 900 0 1 11
0 68
0
0 0 20848 180
2 0V
-7 -16 7 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3512 0 0
2
5.89911e-315 5.40342e-315
0
13 Logic Switch~
5 1889 417 0 1 11
0 92
0
0 0 20848 180
2 0V
-7 -16 7 -8
3 V36
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9912 0 0
2
43746 3
0
13 Logic Switch~
5 1645 108 0 10 11
0 56 0 0 0 0 0 0 0 0
1
0
0 0 20848 180
2 5V
-7 -16 7 -8
3 V31
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3212 0 0
2
43746 4
0
13 Logic Switch~
5 222 1308 0 1 11
0 58
0
0 0 20848 90
2 0V
11 -5 25 3
3 V30
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8247 0 0
2
43746 5
0
13 Logic Switch~
5 195 1128 0 1 11
0 91
0
0 0 20848 90
2 0V
11 -5 25 3
3 V29
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3947 0 0
2
43746 6
0
13 Logic Switch~
5 142 768 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
3 V27
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4251 0 0
2
43746 7
0
13 Logic Switch~
5 35 303 0 1 11
0 137
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -2 0
1 V
938 0 0
2
43746 8
0
13 Logic Switch~
5 626 571 0 1 11
0 93
0
0 0 20848 782
2 0V
-6 -21 8 -13
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
43746 9
0
13 Logic Switch~
5 248 262 0 1 11
0 130
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7643 0 0
2
5.89911e-315 5.4086e-315
0
13 Logic Switch~
5 722 2149 0 10 11
0 138 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
54 68 68 76
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
3236 0 0
2
5.89911e-315 5.41378e-315
0
13 Logic Switch~
5 1057 1528 0 10 11
0 125 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3903 0 0
2
5.89911e-315 5.41896e-315
0
13 Logic Switch~
5 89 67 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3968 0 0
2
5.89911e-315 5.42414e-315
0
13 Logic Switch~
5 433 523 0 1 11
0 103
0
0 0 20848 90
2 0V
-6 15 8 23
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3106 0 0
2
5.89911e-315 5.42933e-315
0
13 Logic Switch~
5 461 523 0 1 11
0 102
0
0 0 20848 90
2 0V
-6 15 8 23
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3223 0 0
2
5.89911e-315 5.43192e-315
0
13 Logic Switch~
5 404 523 0 1 11
0 104
0
0 0 20848 90
2 0V
-6 15 8 23
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6341 0 0
2
5.89911e-315 5.43451e-315
0
13 Logic Switch~
5 373 523 0 1 11
0 105
0
0 0 20848 90
2 0V
-6 15 8 23
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4627 0 0
2
5.89911e-315 5.4371e-315
0
13 Logic Switch~
5 681 459 0 10 11
0 136 0 0 0 0 0 0 0 0
1
0
0 0 20848 512
2 5V
-7 -16 7 -8
2 V5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6952 0 0
2
5.89911e-315 5.43969e-315
0
13 Logic Switch~
5 511 910 0 1 11
0 113
0
0 0 20848 90
2 0V
-6 15 8 23
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3974 0 0
2
5.89911e-315 5.44228e-315
0
13 Logic Switch~
5 539 911 0 1 11
0 112
0
0 0 20848 90
2 0V
-6 15 8 23
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4630 0 0
2
5.89911e-315 5.44487e-315
0
13 Logic Switch~
5 483 910 0 1 11
0 114
0
0 0 20848 90
2 0V
-6 15 8 23
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5705 0 0
2
5.89911e-315 5.44746e-315
0
13 Logic Switch~
5 451 910 0 1 11
0 115
0
0 0 20848 90
2 0V
-6 15 8 23
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8423 0 0
2
5.89911e-315 5.45005e-315
0
13 Logic Switch~
5 611 932 0 10 11
0 135 0 0 0 0 0 0 0 0
1
0
0 0 20848 602
2 5V
11 -5 25 3
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6486 0 0
2
5.89911e-315 5.45264e-315
0
14 Logic Display~
6 1460 658 0 1 2
10 16
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L45
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3367 0 0
2
43746 0
0
14 Logic Display~
6 1451 636 0 1 2
10 17
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L44
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7389 0 0
2
43746 0
0
14 Logic Display~
6 1450 615 0 1 2
10 124
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L43
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6782 0 0
2
43746 0
0
14 Logic Display~
6 1450 599 0 1 2
10 18
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L42
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5728 0 0
2
43746 0
0
14 Logic Display~
6 1530 501 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L41
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6119 0 0
2
43746 0
0
9 Inverter~
13 2336 2200 0 2 22
0 22 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U27A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
3241 0 0
2
43746 0
0
9 Inverter~
13 2518 2693 0 2 22
0 23 11
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U26F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
3835 0 0
2
43746 10
0
7 Ground~
168 1750 372 0 1 3
0 2
0
0 0 53360 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7478 0 0
2
5.89911e-315 5.45523e-315
0
14 Logic Display~
6 1055 1945 0 1 2
10 27
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L22
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3979 0 0
2
5.89911e-315 5.45782e-315
0
14 Logic Display~
6 1053 1901 0 1 2
10 29
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L20
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6285 0 0
2
5.89911e-315 5.46041e-315
0
14 Logic Display~
6 1052 1858 0 1 2
10 24
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L19
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4935 0 0
2
5.89911e-315 5.463e-315
0
14 Logic Display~
6 1052 1833 0 1 2
10 28
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L18
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7650 0 0
2
5.89911e-315 5.46559e-315
0
14 Logic Display~
6 1050 1802 0 1 2
10 30
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L17
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9836 0 0
2
5.89911e-315 5.46818e-315
0
14 Logic Display~
6 1040 1772 0 1 2
10 31
0
0 0 53872 270
6 100MEG
3 -16 45 -8
3 L16
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3988 0 0
2
5.89911e-315 5.47077e-315
0
9 Inverter~
13 991 1949 0 2 22
0 32 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
492 0 0
2
5.89911e-315 5.47207e-315
0
9 Inverter~
13 992 1905 0 2 22
0 33 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
5338 0 0
2
5.89911e-315 5.47336e-315
0
9 Inverter~
13 1002 1861 0 2 22
0 34 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
8324 0 0
2
5.89911e-315 5.47466e-315
0
9 Inverter~
13 1001 1836 0 2 22
0 35 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
9550 0 0
2
5.89911e-315 5.47595e-315
0
9 Inverter~
13 962 1805 0 2 22
0 36 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U26A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
6380 0 0
2
5.89911e-315 5.47725e-315
0
9 Inverter~
13 958 1775 0 2 22
0 37 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U21F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
7942 0 0
2
5.89911e-315 5.47854e-315
0
14 Logic Display~
6 2489 2718 0 1 2
10 23
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L40
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
789 0 0
2
5.89911e-315 5.47984e-315
0
14 Logic Display~
6 2299 2688 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L39
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9884 0 0
2
5.89911e-315 5.48113e-315
0
14 Logic Display~
6 2398 2691 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L38
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6253 0 0
2
5.89911e-315 5.48243e-315
0
14 Logic Display~
6 2372 2686 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L37
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7409 0 0
2
5.89911e-315 5.48372e-315
0
14 Logic Display~
6 2431 2691 0 1 2
10 23
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L36
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3540 0 0
2
5.89911e-315 5.48502e-315
0
14 Logic Display~
6 2338 2688 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L35
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3103 0 0
2
5.89911e-315 5.48631e-315
0
14 Logic Display~
6 2269 2691 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L34
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3548 0 0
2
5.89911e-315 5.48761e-315
0
14 Logic Display~
6 2239 2691 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L33
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9961 0 0
2
5.89911e-315 5.4889e-315
0
14 Logic Display~
6 2158 2695 0 1 2
10 22
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L32
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8521 0 0
2
5.89911e-315 5.4902e-315
0
14 Logic Display~
6 2072 2700 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L31
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5296 0 0
2
5.89911e-315 5.49149e-315
0
14 Logic Display~
6 1968 2698 0 1 2
10 19
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L30
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5398 0 0
2
5.89911e-315 5.49279e-315
0
14 Logic Display~
6 1838 2696 0 1 2
10 14
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L29
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7935 0 0
2
5.89911e-315 5.49408e-315
0
14 Logic Display~
6 1690 2692 0 1 2
10 4
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L28
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
356 0 0
2
5.89911e-315 5.49538e-315
0
14 Logic Display~
6 1494 2706 0 1 2
10 13
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L27
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4629 0 0
2
5.89911e-315 5.49667e-315
0
14 Logic Display~
6 1358 2722 0 1 2
10 15
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L26
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
2
5.89911e-315 5.49797e-315
0
14 Logic Display~
6 1259 2576 0 1 2
10 10
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L25
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5713 0 0
2
5.89911e-315 5.49926e-315
0
14 Logic Display~
6 1163 2508 0 1 2
10 12
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L24
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6618 0 0
2
5.89911e-315 5.50056e-315
0
14 Logic Display~
6 1099 2747 0 1 2
10 9
0
0 0 53872 180
6 100MEG
3 -16 45 -8
3 L23
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3714 0 0
2
5.89911e-315 5.50185e-315
0
8 2-In OR~
219 2140 2543 0 3 22
0 22 39 5
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U23B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
9116 0 0
2
5.89911e-315 5.50315e-315
0
9 2-In AND~
219 2094 2160 0 3 22
0 27 26 22
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U25B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
7960 0 0
2
5.89911e-315 5.50444e-315
0
9 Inverter~
13 2061 2553 0 2 22
0 39 19
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U21E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
3886 0 0
2
5.89911e-315 5.50574e-315
0
9 Inverter~
13 1921 2546 0 2 22
0 40 14
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U21D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
3299 0 0
2
5.89911e-315 5.50703e-315
0
9 2-In AND~
219 2065 2478 0 3 22
0 26 28 39
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U25A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9107 0 0
2
5.89911e-315 5.50833e-315
0
8 2-In OR~
219 1923 2497 0 3 22
0 41 23 40
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U23A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
6556 0 0
2
5.89911e-315 5.50963e-315
0
9 2-In AND~
219 1910 2393 0 3 22
0 29 26 23
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U19B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3205 0 0
2
5.89911e-315 5.51092e-315
0
9 Inverter~
13 1689 2581 0 2 22
0 42 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U21C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
7255 0 0
2
5.89911e-315 5.51222e-315
0
8 2-In OR~
219 1689 2533 0 3 22
0 43 25 42
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U20D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8613 0 0
2
5.89911e-315 5.51286e-315
0
8 2-In OR~
219 1721 2456 0 3 22
0 6 7 43
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U20C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
7832 0 0
2
5.89911e-315 5.51351e-315
0
9 2-In AND~
219 1781 2366 0 3 22
0 26 24 6
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U24D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8937 0 0
2
5.89911e-315 5.51416e-315
0
9 2-In AND~
219 1674 2344 0 3 22
0 26 30 7
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U24C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
556 0 0
2
5.89911e-315 5.51481e-315
0
9 Inverter~
13 1489 2319 0 2 22
0 44 13
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U21B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
6981 0 0
2
5.89911e-315 5.51545e-315
0
8 2-In OR~
219 1488 2273 0 3 22
0 25 10 44
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U20B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8701 0 0
2
5.89911e-315 5.5161e-315
0
9 2-In AND~
219 1497 2197 0 3 22
0 45 31 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U24B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5540 0 0
2
5.89911e-315 5.51675e-315
0
9 Inverter~
13 1353 2243 0 2 22
0 10 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U21A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
8365 0 0
2
5.89911e-315 5.5174e-315
0
9 Inverter~
13 1139 2264 0 2 22
0 46 12
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U18F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
5209 0 0
2
5.89911e-315 5.51804e-315
0
8 2-In OR~
219 1139 2177 0 3 22
0 41 9 46
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U20A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3297 0 0
2
5.89911e-315 5.51869e-315
0
9 2-In AND~
219 1159 2108 0 3 22
0 31 26 41
0
0 0 624 270
5 74F08
-18 -24 17 -16
4 U19A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9904 0 0
2
5.89911e-315 5.51934e-315
0
9 Inverter~
13 315 1735 0 2 22
0 139 140
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U18C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 3 2 0
1 U
6918 0 0
2
5.89911e-315 5.51999e-315
0
7 Ground~
168 588 1927 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7751 0 0
2
5.89911e-315 5.52063e-315
0
7 74LS154
95 818 1901 0 22 45
0 2 2 48 49 50 47 141 142 143
144 145 146 147 148 149 150 32 33 34
35 36 37
0
0 0 4848 692
7 74LS154
-24 -87 25 -79
3 U15
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 512 1 0 0 0
1 U
9907 0 0
2
43746 11
0
9 Inverter~
13 392 868 0 2 22
0 151 20
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U22D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 4 1 0
1 U
6628 0 0
2
43746 12
0
14 Logic Display~
6 737 50 0 1 2
10 124
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4914 0 0
2
43746 13
0
12 SPST Switch~
165 460 706 0 2 11
0 54 13
0
0 0 4208 0
0
2 S1
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
635 0 0
2
43746 14
0
14 Logic Display~
6 1622 974 0 1 2
10 152
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3606 0 0
2
43746 15
0
7 Ground~
168 1496 552 0 1 3
0 2
0
0 0 53360 692
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
8769 0 0
2
5.89911e-315 5.52128e-315
0
9 Inverter~
13 417 781 0 2 22
0 59 153
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U22C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 3 1 0
1 U
3887 0 0
2
5.89911e-315 5.52193e-315
0
9 Inverter~
13 303 810 0 2 22
0 154 60
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U22B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 2 1 0
1 U
4266 0 0
2
5.89911e-315 5.52258e-315
0
9 2-In AND~
219 367 801 0 3 22
0 61 60 59
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U24A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3389 0 0
2
5.89911e-315 5.52322e-315
0
7 Ground~
168 1453 759 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
8108 0 0
2
43746 16
0
7 74LS157
122 1533 748 0 14 29
0 6 80 76 78 16 77 17 79 18
75 70 71 73 72
0
0 0 4336 270
7 74LS157
-24 -60 25 -52
3 U35
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3301 0 0
2
43746 17
0
7 Ground~
168 1895 570 0 1 3
0 2
0
0 0 53360 180
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3739 0 0
2
43746 18
0
7 74LS173
129 1836 642 0 14 29
0 2 55 155 124 67 68 69 62 2
2 79 77 78 80
0
0 0 4336 0
7 74LS173
-24 -51 25 -43
3 U34
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
4610 0 0
2
43746 19
0
14 Logic Display~
6 1013 1332 0 1 2
10 81
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L319
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7104 0 0
2
5.89911e-315 5.52387e-315
0
14 Logic Display~
6 984 1332 0 1 2
10 82
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L318
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5233 0 0
2
5.89911e-315 5.52452e-315
0
14 Logic Display~
6 954 1332 0 1 2
10 83
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L317
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
345 0 0
2
5.89911e-315 5.52517e-315
0
14 Logic Display~
6 924 1332 0 1 2
10 61
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L316
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4311 0 0
2
5.89911e-315 5.52581e-315
0
14 Logic Display~
6 867 1332 0 1 2
10 85
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L315
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3959 0 0
2
5.89911e-315 5.52646e-315
0
14 Logic Display~
6 836 1332 0 1 2
10 86
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L314
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9550 0 0
2
5.89911e-315 5.52711e-315
0
14 Logic Display~
6 804 1331 0 1 2
10 87
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L313
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4183 0 0
2
5.89911e-315 5.52776e-315
0
14 Logic Display~
6 772 1331 0 1 2
10 88
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L312
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7662 0 0
2
5.89911e-315 5.52841e-315
0
14 Logic Display~
6 772 962 0 1 2
10 88
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L311
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6373 0 0
2
5.89911e-315 5.52905e-315
0
14 Logic Display~
6 804 962 0 1 2
10 87
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L310
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
76 0 0
2
5.89911e-315 5.5297e-315
0
14 Logic Display~
6 836 962 0 1 2
10 86
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L309
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4168 0 0
2
5.89911e-315 5.53035e-315
0
14 Logic Display~
6 867 962 0 1 2
10 85
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L308
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9490 0 0
2
5.89911e-315 5.531e-315
0
14 Logic Display~
6 924 962 0 1 2
10 61
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L307
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3202 0 0
2
5.89911e-315 5.53164e-315
0
14 Logic Display~
6 954 962 0 1 2
10 83
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L306
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5212 0 0
2
5.89911e-315 5.53229e-315
0
14 Logic Display~
6 984 962 0 1 2
10 82
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L305
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5341 0 0
2
5.89911e-315 5.53294e-315
0
14 Logic Display~
6 1013 961 0 1 2
10 81
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L304
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3516 0 0
2
5.89911e-315 5.53359e-315
0
14 Logic Display~
6 772 586 0 1 2
10 88
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L303
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6823 0 0
2
5.89911e-315 5.53423e-315
0
14 Logic Display~
6 804 586 0 1 2
10 87
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L302
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3532 0 0
2
5.89911e-315 5.53488e-315
0
14 Logic Display~
6 836 585 0 1 2
10 86
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L301
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3978 0 0
2
5.89911e-315 5.53553e-315
0
14 Logic Display~
6 867 585 0 1 2
10 85
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L300
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4691 0 0
2
5.89911e-315 5.53618e-315
0
14 Logic Display~
6 924 586 0 1 2
10 61
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L299
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5392 0 0
2
5.89911e-315 5.53682e-315
0
14 Logic Display~
6 954 586 0 1 2
10 83
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L298
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3264 0 0
2
5.89911e-315 5.53747e-315
0
14 Logic Display~
6 984 586 0 1 2
10 82
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L297
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7602 0 0
2
5.89911e-315 5.53812e-315
0
14 Logic Display~
6 1013 586 0 1 2
10 81
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L296
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4228 0 0
2
5.89911e-315 5.53877e-315
0
14 Logic Display~
6 612 274 0 1 2
10 81
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L287
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8797 0 0
2
5.89911e-315 5.53941e-315
0
14 Logic Display~
6 612 256 0 1 2
10 82
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L286
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5117 0 0
2
5.89911e-315 5.54006e-315
0
14 Logic Display~
6 612 238 0 1 2
10 83
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L285
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5387 0 0
2
5.89911e-315 5.54071e-315
0
14 Logic Display~
6 612 220 0 1 2
10 61
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L284
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6535 0 0
2
5.89911e-315 5.54136e-315
0
14 Logic Display~
6 488 274 0 1 2
10 94
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L283
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8927 0 0
2
5.89911e-315 5.542e-315
0
14 Logic Display~
6 488 256 0 1 2
10 95
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L282
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5209 0 0
2
5.89911e-315 5.54265e-315
0
14 Logic Display~
6 488 238 0 1 2
10 96
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L281
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9271 0 0
2
5.89911e-315 5.5433e-315
0
14 Logic Display~
6 488 220 0 1 2
10 97
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L280
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4455 0 0
2
5.89911e-315 5.54395e-315
0
14 Logic Display~
6 335 277 0 1 2
10 81
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L279
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8623 0 0
2
5.89911e-315 5.54459e-315
0
14 Logic Display~
6 321 267 0 1 2
10 82
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L278
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7340 0 0
2
5.89911e-315 5.54524e-315
0
14 Logic Display~
6 304 259 0 1 2
10 83
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L277
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6167 0 0
2
5.89911e-315 5.54589e-315
0
14 Logic Display~
6 290 250 0 1 2
10 61
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L276
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7993 0 0
2
5.89911e-315 5.54654e-315
0
14 Logic Display~
6 722 345 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L275
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3144 0 0
2
5.89911e-315 5.54719e-315
0
14 Logic Display~
6 700 327 0 1 2
10 82
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L274
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3180 0 0
2
5.89911e-315 5.54783e-315
0
14 Logic Display~
6 673 308 0 1 2
10 83
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L273
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7665 0 0
2
5.89911e-315 5.54848e-315
0
14 Logic Display~
6 649 292 0 1 2
10 61
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L272
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7757 0 0
2
5.89911e-315 5.54913e-315
0
14 Logic Display~
6 617 446 0 1 2
10 98
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L271
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4319 0 0
2
5.89911e-315 5.54978e-315
0
14 Logic Display~
6 599 437 0 1 2
10 99
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L270
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7554 0 0
2
5.89911e-315 5.55042e-315
0
14 Logic Display~
6 581 427 0 1 2
10 100
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L269
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
453 0 0
2
5.89911e-315 5.55107e-315
0
14 Logic Display~
6 563 420 0 1 2
10 101
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L268
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9688 0 0
2
5.89911e-315 5.55172e-315
0
14 Logic Display~
6 462 492 0 1 2
10 102
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L267
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8216 0 0
2
5.89911e-315 5.55237e-315
0
14 Logic Display~
6 434 492 0 1 2
10 103
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L266
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3830 0 0
2
5.89911e-315 5.55301e-315
0
14 Logic Display~
6 405 492 0 1 2
10 104
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L265
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3215 0 0
2
5.89911e-315 5.55366e-315
0
14 Logic Display~
6 374 492 0 1 2
10 105
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L264
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3894 0 0
2
5.89911e-315 5.55398e-315
0
14 Logic Display~
6 608 635 0 1 2
10 106
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L263
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3490 0 0
2
5.89911e-315 5.55431e-315
0
14 Logic Display~
6 590 635 0 1 2
10 107
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L262
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5596 0 0
2
5.89911e-315 5.55463e-315
0
14 Logic Display~
6 572 635 0 1 2
10 108
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L261
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3848 0 0
2
5.89911e-315 5.55496e-315
0
14 Logic Display~
6 554 635 0 1 2
10 109
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L260
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6792 0 0
2
5.89911e-315 5.55528e-315
0
14 Logic Display~
6 745 707 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L259
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
756 0 0
2
5.89911e-315 5.5556e-315
0
14 Logic Display~
6 745 698 0 1 2
10 82
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L258
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6249 0 0
2
5.89911e-315 5.55593e-315
0
14 Logic Display~
6 745 689 0 1 2
10 83
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L257
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3967 0 0
2
5.89911e-315 5.55625e-315
0
14 Logic Display~
6 745 680 0 1 2
10 61
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L256
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.89911e-315 5.55657e-315
0
14 Logic Display~
6 745 671 0 1 2
10 85
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L255
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3435 0 0
2
5.89911e-315 5.5569e-315
0
14 Logic Display~
6 745 662 0 1 2
10 86
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L254
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7674 0 0
2
5.89911e-315 5.55722e-315
0
14 Logic Display~
6 745 653 0 1 2
10 87
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L253
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3516 0 0
2
5.89911e-315 5.55755e-315
0
14 Logic Display~
6 745 644 0 1 2
10 88
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L252
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6731 0 0
2
5.89911e-315 5.55787e-315
0
14 Logic Display~
6 725 738 0 1 2
10 89
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L251
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3620 0 0
2
5.89911e-315 5.55819e-315
0
14 Logic Display~
6 707 738 0 1 2
10 90
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L250
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
5.89911e-315 5.55852e-315
0
14 Logic Display~
6 671 738 0 1 2
10 110
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L248
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3480 0 0
2
5.89911e-315 5.55884e-315
0
14 Logic Display~
6 689 737 0 1 2
10 111
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L249
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8526 0 0
2
5.89911e-315 5.55917e-315
0
14 Logic Display~
6 734 881 0 1 2
10 81
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L247
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7437 0 0
2
5.89911e-315 5.55949e-315
0
14 Logic Display~
6 716 881 0 1 2
10 82
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L246
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8275 0 0
2
5.89911e-315 5.55981e-315
0
14 Logic Display~
6 698 882 0 1 2
10 83
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L245
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6488 0 0
2
5.89911e-315 5.56014e-315
0
14 Logic Display~
6 680 882 0 1 2
10 61
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L244
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3483 0 0
2
5.89911e-315 5.56046e-315
0
14 Logic Display~
6 540 874 0 1 2
10 112
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L243
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4998 0 0
2
5.89911e-315 5.56078e-315
0
14 Logic Display~
6 512 874 0 1 2
10 113
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L242
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5846 0 0
2
5.89911e-315 5.56111e-315
0
14 Logic Display~
6 484 874 0 1 2
10 114
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L241
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3129 0 0
2
5.89911e-315 5.56143e-315
0
14 Logic Display~
6 452 874 0 1 2
10 115
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L240
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4249 0 0
2
5.89911e-315 5.56176e-315
0
14 Logic Display~
6 705 1157 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L239
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9669 0 0
2
5.89911e-315 5.56208e-315
0
14 Logic Display~
6 684 1148 0 1 2
10 82
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L238
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5459 0 0
2
5.89911e-315 5.5624e-315
0
14 Logic Display~
6 665 1139 0 1 2
10 83
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L237
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3156 0 0
2
5.89911e-315 5.56273e-315
0
14 Logic Display~
6 646 1130 0 1 2
10 61
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L236
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4876 0 0
2
5.89911e-315 5.56305e-315
0
14 Logic Display~
6 471 1273 0 1 2
10 85
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L235
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3723 0 0
2
5.89911e-315 5.56337e-315
0
14 Logic Display~
6 457 1263 0 1 2
10 86
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L234
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3827 0 0
2
5.89911e-315 5.5637e-315
0
14 Logic Display~
6 446 1254 0 1 2
10 87
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L233
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
70 0 0
2
5.89911e-315 5.56402e-315
0
14 Logic Display~
6 435 1244 0 1 2
10 88
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L232
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4465 0 0
2
5.89911e-315 5.56435e-315
0
14 Logic Display~
6 510 1357 0 1 2
10 47
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L231
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8698 0 0
2
5.89911e-315 5.56467e-315
0
14 Logic Display~
6 519 1336 0 1 2
10 50
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L230
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4766 0 0
2
5.89911e-315 5.56499e-315
0
14 Logic Display~
6 528 1315 0 1 2
10 49
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L229
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8576 0 0
2
5.89911e-315 5.56532e-315
0
14 Logic Display~
6 538 1299 0 1 2
10 48
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L228
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
5.89911e-315 5.56564e-315
0
14 Logic Display~
6 757 1110 0 1 2
10 81
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L227
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9662 0 0
2
5.89911e-315 5.56596e-315
0
14 Logic Display~
6 750 1101 0 1 2
10 82
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L226
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3374 0 0
2
5.89911e-315 5.56629e-315
0
14 Logic Display~
6 739 1092 0 1 2
10 83
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L225
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4396 0 0
2
5.89911e-315 5.56661e-315
0
14 Logic Display~
6 726 1083 0 1 2
10 61
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L224
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5842 0 0
2
5.89911e-315 5.56694e-315
0
14 Logic Display~
6 1046 544 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L222
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6972 0 0
2
5.89911e-315 5.56726e-315
0
14 Logic Display~
6 1046 526 0 1 2
10 82
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L221
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3913 0 0
2
5.89911e-315 5.56758e-315
0
14 Logic Display~
6 1046 508 0 1 2
10 83
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L220
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4772 0 0
2
5.89911e-315 5.56791e-315
0
14 Logic Display~
6 1046 490 0 1 2
10 61
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L219
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8158 0 0
2
5.89911e-315 5.56823e-315
0
14 Logic Display~
6 1046 341 0 1 2
10 81
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L218
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5328 0 0
2
5.89911e-315 5.56856e-315
0
14 Logic Display~
6 1046 323 0 1 2
10 82
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L217
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3402 0 0
2
5.89911e-315 5.56888e-315
0
14 Logic Display~
6 1046 305 0 1 2
10 83
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L216
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9932 0 0
2
5.89911e-315 5.5692e-315
0
14 Logic Display~
6 1046 287 0 1 2
10 61
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L215
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3452 0 0
2
5.89911e-315 5.56953e-315
0
14 Logic Display~
6 1170 342 0 1 2
10 116
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L214
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9735 0 0
2
5.89911e-315 5.56985e-315
0
14 Logic Display~
6 1170 323 0 1 2
10 117
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L213
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
493 0 0
2
5.89911e-315 5.57017e-315
0
14 Logic Display~
6 1170 305 0 1 2
10 118
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L212
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4627 0 0
2
5.89911e-315 5.5705e-315
0
14 Logic Display~
6 1169 287 0 1 2
10 119
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L211
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3860 0 0
2
5.89911e-315 5.57082e-315
0
14 Logic Display~
6 1146 544 0 1 2
10 120
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L210
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5167 0 0
2
5.89911e-315 5.57115e-315
0
14 Logic Display~
6 1146 526 0 1 2
10 121
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L209
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4856 0 0
2
5.89911e-315 5.57147e-315
0
14 Logic Display~
6 1146 508 0 1 2
10 122
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L208
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3839 0 0
2
5.89911e-315 5.57179e-315
0
14 Logic Display~
6 1146 490 0 1 2
10 123
0
0 0 53360 782
6 100MEG
3 -16 45 -8
4 L207
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8865 0 0
2
5.89911e-315 5.57212e-315
0
14 Logic Display~
6 1349 427 0 1 2
10 116
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L201
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7317 0 0
2
5.89911e-315 5.57244e-315
0
14 Logic Display~
6 1335 427 0 1 2
10 117
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L200
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
372 0 0
2
5.89911e-315 5.57276e-315
0
14 Logic Display~
6 1321 427 0 1 2
10 118
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L199
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7592 0 0
2
5.89911e-315 5.57309e-315
0
14 Logic Display~
6 1308 427 0 1 2
10 119
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L198
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3434 0 0
2
5.89911e-315 5.57341e-315
0
14 Logic Display~
6 1349 245 0 1 2
10 116
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L197
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
367 0 0
2
5.89911e-315 5.57374e-315
0
14 Logic Display~
6 1335 245 0 1 2
10 117
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L196
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
35 0 0
2
5.89911e-315 5.57406e-315
0
14 Logic Display~
6 1321 245 0 1 2
10 118
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L195
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4461 0 0
2
5.89911e-315 5.57438e-315
0
14 Logic Display~
6 1308 245 0 1 2
10 119
0
0 0 53360 692
6 100MEG
3 -16 45 -8
4 L194
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7455 0 0
2
5.89911e-315 5.57471e-315
0
14 Logic Display~
6 1129 930 0 1 2
10 81
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L187
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5237 0 0
2
5.89911e-315 5.57503e-315
0
14 Logic Display~
6 1108 921 0 1 2
10 82
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L186
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5896 0 0
2
5.89911e-315 5.57535e-315
0
14 Logic Display~
6 1085 912 0 1 2
10 83
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L185
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4980 0 0
2
5.89911e-315 5.57568e-315
0
14 Logic Display~
6 1065 902 0 1 2
10 61
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L184
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
367 0 0
2
5.89911e-315 5.576e-315
0
14 Logic Display~
6 1125 221 0 1 2
10 81
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L183
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5653 0 0
2
5.89911e-315 5.57633e-315
0
14 Logic Display~
6 1101 212 0 1 2
10 82
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L182
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4544 0 0
2
5.89911e-315 5.57665e-315
0
14 Logic Display~
6 1076 203 0 1 2
10 83
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L181
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6756 0 0
2
5.89911e-315 5.57697e-315
0
14 Logic Display~
6 1055 194 0 1 2
10 61
0
0 0 53360 602
6 100MEG
3 -16 45 -8
4 L180
-15 -15 13 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6495 0 0
2
5.89911e-315 5.5773e-315
0
12 SPST Switch~
165 741 1470 0 10 11
0 124 124 0 0 0 0 0 0 0
1
0
0 0 4208 0
0
2 S7
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3703 0 0
2
5.89911e-315 5.57762e-315
0
9 Terminal~
194 648 1461 0 1 3
0 124
0
0 0 49520 0
3 CLK
-11 -22 10 -14
3 T21
-11 -32 10 -24
0
4 CLK;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3988 0 0
2
5.89911e-315 5.57795e-315
0
14 Logic Display~
6 2761 3065 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L174
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6270 0 0
2
43746 20
0
14 Logic Display~
6 2732 2978 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L173
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3193 0 0
2
43746 21
0
14 Logic Display~
6 2703 2902 0 1 2
10 156
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L172
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
7594 0 0
2
43746 22
0
14 Logic Display~
6 2671 2820 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L171
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7298 0 0
2
43746 23
0
14 Logic Display~
6 2641 2746 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L170
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3595 0 0
2
43746 24
0
14 Logic Display~
6 2611 2670 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L169
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
464 0 0
2
43746 25
0
14 Logic Display~
6 2581 2598 0 1 2
10 157
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L168
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
8913 0 0
2
43746 26
0
14 Logic Display~
6 2551 2530 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L167
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8648 0 0
2
43746 27
0
14 Logic Display~
6 2522 2448 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L166
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3202 0 0
2
43746 28
0
14 Logic Display~
6 2463 2290 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L164
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5604 0 0
2
43746 29
0
14 Logic Display~
6 2762 2258 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L163
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8890 0 0
2
43746 30
0
14 Logic Display~
6 2731 2236 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L162
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7714 0 0
2
43746 31
0
14 Logic Display~
6 2704 2214 0 1 2
10 158
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L161
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
366 0 0
2
43746 32
0
14 Logic Display~
6 2671 2188 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L160
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8936 0 0
2
43746 33
0
14 Logic Display~
6 2642 2168 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L159
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6354 0 0
2
43746 34
0
14 Logic Display~
6 2612 2140 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L158
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9149 0 0
2
43746 35
0
14 Logic Display~
6 2583 2120 0 1 2
10 159
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L157
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
382 0 0
2
43746 36
0
14 Logic Display~
6 2551 2100 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L156
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3142 0 0
2
43746 37
0
14 Logic Display~
6 2522 2074 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L155
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6989 0 0
2
43746 38
0
14 Logic Display~
6 2463 2018 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L153
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3569 0 0
2
43746 39
0
14 Logic Display~
6 2761 1730 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L152
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4568 0 0
2
43746 40
0
14 Logic Display~
6 2732 1714 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L151
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6294 0 0
2
43746 41
0
14 Logic Display~
6 2670 1678 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L149
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9900 0 0
2
43746 42
0
14 Logic Display~
6 2641 1662 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L148
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6441 0 0
2
43746 43
0
14 Logic Display~
6 2611 1650 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L147
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
780 0 0
2
43746 44
0
14 Logic Display~
6 2581 1634 0 1 2
10 160
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L146
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3797 0 0
2
43746 45
0
14 Logic Display~
6 2551 1618 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L145
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
371 0 0
2
43746 46
0
14 Logic Display~
6 2522 1598 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L144
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6265 0 0
2
43746 47
0
14 Logic Display~
6 2463 1531 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L142
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5116 0 0
2
43746 48
0
14 Logic Display~
6 2463 1531 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L141
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4818 0 0
2
43746 49
0
14 Logic Display~
6 2762 1307 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L140
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3119 0 0
2
43746 50
0
14 Logic Display~
6 2733 1286 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L139
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
656 0 0
2
43746 51
0
14 Logic Display~
6 2671 1251 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L137
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9129 0 0
2
43746 52
0
14 Logic Display~
6 2642 1230 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L136
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8217 0 0
2
43746 53
0
14 Logic Display~
6 2612 1204 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L135
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9758 0 0
2
43746 54
0
14 Logic Display~
6 2583 1190 0 1 2
10 161
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L134
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3132 0 0
2
43746 55
0
14 Logic Display~
6 2551 1170 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L133
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4637 0 0
2
43746 56
0
14 Logic Display~
6 2522 1152 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L132
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3390 0 0
2
43746 57
0
14 Logic Display~
6 2463 1113 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L130
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8561 0 0
2
43746 58
0
14 Logic Display~
6 2761 544 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L129
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6596 0 0
2
43746 59
0
14 Logic Display~
6 2732 520 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L128
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
829 0 0
2
43746 60
0
14 Logic Display~
6 2671 470 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L126
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7394 0 0
2
43746 61
0
14 Logic Display~
6 2641 450 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L125
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6213 0 0
2
43746 62
0
14 Logic Display~
6 2611 548 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L124
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4924 0 0
2
43746 63
0
14 Logic Display~
6 2582 530 0 1 2
10 162
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L123
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
975 0 0
2
43746 64
0
14 Logic Display~
6 2551 519 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L122
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4193 0 0
2
43746 65
0
14 Logic Display~
6 2522 505 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L121
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7871 0 0
2
43746 66
0
14 Logic Display~
6 2761 903 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L120
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7844 0 0
2
43746 67
0
14 Logic Display~
6 2732 882 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L119
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4539 0 0
2
43746 68
0
14 Logic Display~
6 2671 847 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L117
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6378 0 0
2
43746 69
0
14 Logic Display~
6 2641 824 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L116
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
733 0 0
2
43746 70
0
14 Logic Display~
6 2611 798 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L115
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3524 0 0
2
43746 71
0
14 Logic Display~
6 2581 777 0 1 2
10 163
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L114
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
3286 0 0
2
43746 72
0
14 Logic Display~
6 2552 755 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L113
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6414 0 0
2
43746 73
0
14 Logic Display~
6 2522 732 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L112
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
381 0 0
2
43746 74
0
14 Logic Display~
6 27 2738 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L110
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
456 0 0
2
43746 75
0
14 Logic Display~
6 57 2680 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L109
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3688 0 0
2
43746 76
0
14 Logic Display~
6 85 2616 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L108
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3367 0 0
2
43746 77
0
14 Logic Display~
6 113 2552 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L107
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3557 0 0
2
43746 78
0
14 Logic Display~
6 169 2424 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L105
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7241 0 0
2
43746 79
0
14 Logic Display~
6 196 2363 0 1 2
10 14
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L104
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4540 0 0
2
43746 80
0
14 Logic Display~
6 223 2309 0 1 2
10 15
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L103
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4740 0 0
2
43746 81
0
14 Logic Display~
6 224 2044 0 1 2
10 15
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L102
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9311 0 0
2
43746 82
0
14 Logic Display~
6 196 1997 0 1 2
10 14
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L101
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5668 0 0
2
43746 83
0
14 Logic Display~
6 169 1949 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
4 L100
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7265 0 0
2
43746 84
0
14 Logic Display~
6 113 1832 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L98
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7410 0 0
2
43746 85
0
14 Logic Display~
6 86 1776 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L97
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3365 0 0
2
43746 86
0
14 Logic Display~
6 57 1726 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L96
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4709 0 0
2
43746 87
0
14 Logic Display~
6 28 1686 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L95
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9224 0 0
2
43746 88
0
14 Logic Display~
6 223 1432 0 1 2
10 15
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L94
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
43746 89
0
14 Logic Display~
6 196 1376 0 1 2
10 14
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L93
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
372 0 0
2
43746 90
0
14 Logic Display~
6 169 1330 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L92
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3192 0 0
2
43746 91
0
14 Logic Display~
6 115 1248 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L90
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3923 0 0
2
43746 92
0
14 Logic Display~
6 85 1212 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L89
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6312 0 0
2
43746 93
0
14 Logic Display~
6 57 1166 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L88
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3973 0 0
2
43746 94
0
14 Logic Display~
6 28 1122 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L87
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3791 0 0
2
43746 95
0
14 Logic Display~
6 223 1173 0 1 2
10 15
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L86
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5134 0 0
2
43746 96
0
14 Logic Display~
6 196 1008 0 1 2
10 14
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L85
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3564 0 0
2
43746 97
0
14 Logic Display~
6 169 906 0 1 2
10 13
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L84
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9962 0 0
2
43746 98
0
14 Logic Display~
6 114 824 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L82
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4113 0 0
2
43746 99
0
14 Logic Display~
6 86 770 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L81
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4683 0 0
2
43746 100
0
14 Logic Display~
6 57 731 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L80
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6923 0 0
2
43746 101
0
14 Logic Display~
6 28 707 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L79
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8938 0 0
2
43746 102
0
14 Logic Display~
6 114 518 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L78
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
975 0 0
2
43746 103
0
14 Logic Display~
6 57 430 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L76
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9382 0 0
2
43746 104
0
14 Logic Display~
6 28 396 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L75
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3443 0 0
2
43746 105
0
14 Logic Display~
6 532 105 0 1 2
10 9
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L74
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8770 0 0
2
43746 106
0
14 Logic Display~
6 194 104 0 1 2
10 9
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L73
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5396 0 0
2
43746 107
0
14 Logic Display~
6 159 206 0 1 2
10 10
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L72
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6225 0 0
2
43746 108
0
14 Logic Display~
6 193 301 0 1 2
10 12
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L70
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9851 0 0
2
43746 109
0
14 Logic Display~
6 189 641 0 1 2
10 20
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L69
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3954 0 0
2
43746 110
0
14 Logic Display~
6 189 670 0 1 2
10 13
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L68
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7375 0 0
2
43746 111
0
14 Logic Display~
6 1619 810 0 1 2
10 84
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L67
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
699 0 0
2
43746 112
0
14 Logic Display~
6 1611 574 0 1 2
10 164
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L66
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
6991 0 0
2
43746 113
0
14 Logic Display~
6 1729 473 0 1 2
10 6
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L65
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7573 0 0
2
43746 114
0
14 Logic Display~
6 1692 464 0 1 2
10 7
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L64
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8781 0 0
2
43746 115
0
14 Logic Display~
6 1650 455 0 1 2
10 7
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L63
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9995 0 0
2
43746 116
0
14 Logic Display~
6 1610 445 0 1 2
10 6
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L62
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6952 0 0
2
43746 117
0
14 Logic Display~
6 1610 397 0 1 2
10 7
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L61
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9357 0 0
2
43746 118
0
14 Logic Display~
6 1610 377 0 1 2
10 6
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L60
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5834 0 0
2
43746 119
0
14 Logic Display~
6 1610 358 0 1 2
10 2
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L59
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3722 0 0
2
43746 120
0
14 Logic Display~
6 1607 266 0 1 2
10 5
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L58
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8504 0 0
2
43746 121
0
14 Logic Display~
6 1602 105 0 1 2
10 4
0
0 0 53360 90
6 100MEG
3 -16 45 -8
3 L57
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8638 0 0
2
43746 122
0
7 Pulser~
4 834 1518 0 11 12
0 38 165 124 166 0 0 10 10 -1
7 1
0
0 0 4144 0
0
3 V14
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
389 0 0
2
5.89911e-315 5.57827e-315
0
9 Terminal~
194 2761 3121 0 1 3
0 4
0
0 0 49520 180
5 LaBAR
6 -7 41 1
3 T19
-11 -32 10 -24
0
6 LaBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7306 0 0
2
5.89911e-315 5.57859e-315
0
9 Terminal~
194 2732 3039 0 1 3
0 5
0
0 0 49520 180
2 Ea
-5 -1 9 7
3 T18
-10 -32 11 -24
0
3 Ea;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
434 0 0
2
5.89911e-315 5.57892e-315
0
9 Terminal~
194 2704 2956 0 1 3
0 0
0
0 0 49520 180
2 Eu
-5 1 9 9
3 T17
-10 -32 11 -24
0
3 Eu;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
7417 0 0
2
5.89911e-315 5.57924e-315
0
9 Terminal~
194 2671 2872 0 1 3
0 6
0
0 0 49520 180
1 M
-3 -1 4 7
3 T16
-11 -32 10 -24
0
2 M;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
320 0 0
2
5.89911e-315 5.57956e-315
0
9 Terminal~
194 2641 2800 0 1 3
0 7
0
0 0 49520 180
3 Cin
-9 -1 12 7
3 T15
-11 -32 10 -24
0
4 Cin;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7907 0 0
2
5.89911e-315 5.57989e-315
0
9 Terminal~
194 2611 2731 0 1 3
0 6
0
0 0 49520 180
2 S3
-6 -2 8 6
3 T14
-10 -32 11 -24
0
3 S3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7378 0 0
2
5.89911e-315 5.58021e-315
0
9 Terminal~
194 2582 2652 0 1 3
0 0
0
0 0 49520 180
2 S2
-5 0 9 8
3 T13
-10 -32 11 -24
0
3 S2;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
7918 0 0
2
5.89911e-315 5.58054e-315
0
9 Terminal~
194 2576 2776 0 1 3
0 7
0
0 0 49520 180
2 S1
-6 -1 8 7
3 T12
-10 -32 11 -24
0
3 S1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6109 0 0
2
5.89911e-315 5.58086e-315
0
9 Terminal~
194 2522 2497 0 1 3
0 6
0
0 0 49520 180
2 S0
7 -7 21 1
3 T11
-10 -32 11 -24
0
3 S0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3630 0 0
2
5.89911e-315 5.58118e-315
0
9 Terminal~
194 2464 2337 0 1 3
0 8
0
0 0 49520 692
5 LoBAR
-16 -1 19 7
2 T9
-8 -32 6 -24
0
6 LoBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3956 0 0
2
5.89911e-315 5.58151e-315
0
9 Terminal~
194 28 2783 0 1 3
0 9
0
0 0 49520 180
2 Ep
-7 0 7 8
2 T8
-7 -32 7 -24
0
3 Ep;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
350 0 0
2
5.89911e-315 5.58183e-315
0
9 Terminal~
194 57 2720 0 1 3
0 10
0
0 0 49520 180
2 Cp
-6 0 8 8
2 T7
-7 -32 7 -24
0
3 Cp;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
326 0 0
2
5.89911e-315 5.58215e-315
0
9 Terminal~
194 86 2662 0 1 3
0 11
0
0 0 49520 180
5 LpBAR
-16 -1 19 7
2 T6
-7 -32 7 -24
0
6 LpBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9825 0 0
2
5.89911e-315 5.58248e-315
0
9 Terminal~
194 114 2600 0 1 3
0 12
0
0 0 49520 180
5 LmBAR
-16 -1 19 7
2 T5
-8 -32 6 -24
0
6 LmBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8211 0 0
2
5.89911e-315 5.5828e-315
0
9 Terminal~
194 169 2470 0 1 3
0 13
0
0 0 49520 180
5 CEbar
-17 -1 18 7
2 T3
-8 -32 6 -24
0
6 CEbar;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7360 0 0
2
5.89911e-315 5.58313e-315
0
9 Terminal~
194 226 2473 0 1 3
0 14
0
0 0 49520 180
5 EiBAR
-16 -1 19 7
2 T2
-8 -32 6 -24
0
6 EiBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7114 0 0
2
5.89911e-315 5.58345e-315
0
9 Terminal~
194 223 2354 0 1 3
0 15
0
0 0 49520 180
5 LiBAR
-17 -1 18 7
2 T1
-7 -32 7 -24
0
6 LiBAR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3107 0 0
2
5.89911e-315 5.58377e-315
0
14 Logic Display~
6 927 1623 0 1 2
10 9
0
0 0 53360 270
6 100MEG
3 -16 45 -8
3 L10
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8732 0 0
2
5.89911e-315 5.5841e-315
0
14 Logic Display~
6 927 1650 0 1 2
10 10
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L9
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6705 0 0
2
5.89911e-315 5.58442e-315
0
14 Logic Display~
6 927 1680 0 1 2
10 26
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L8
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7374 0 0
2
5.89911e-315 5.58474e-315
0
14 Logic Display~
6 927 1708 0 1 2
10 45
0
0 0 53360 270
6 100MEG
3 -16 45 -8
2 L7
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6457 0 0
2
5.89911e-315 5.58507e-315
0
14 Logic Display~
6 2288 1709 0 1 2
10 45
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L14
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3501 0 0
2
43746 123
0
14 Logic Display~
6 2287 1681 0 1 2
10 26
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L13
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9597 0 0
2
43746 124
0
14 Logic Display~
6 2287 1651 0 1 2
10 10
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L12
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9950 0 0
2
43746 125
0
14 Logic Display~
6 2287 1624 0 1 2
10 9
0
0 0 53360 602
6 100MEG
3 -16 45 -8
3 L11
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3239 0 0
2
43746 126
0
14 Logic Display~
6 1025 1434 0 1 2
10 124
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7621 0 0
2
5.89911e-315 5.58539e-315
0
7 74LS107
112 1439 1476 0 12 25
0 128 45 124 125 9 127 124 125 127
9 10 126
0
0 0 4336 0
7 74LS107
-24 -51 25 -43
3 U17
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 4 12 13 8 11 9 10 3
2 5 6 1 4 12 13 8 11 9
10 3 2 5 6 0
65 0 0 0 1 1 0 0
1 U
8673 0 0
2
5.89911e-315 5.58572e-315
0
7 74LS107
112 1214 1479 0 12 25
0 10 126 124 125 26 129 124 125 26
129 45 128
0
0 0 4336 0
7 74LS107
-24 -51 25 -43
3 U16
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 4 12 13 8 11 9 10 3
2 5 6 1 4 12 13 8 11 9
10 3 2 5 6 0
65 0 0 0 1 0 0 0
1 U
9712 0 0
2
5.89911e-315 5.58604e-315
0
14 Logic Display~
6 221 32 0 1 2
10 124
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3900 0 0
2
5.89911e-315 5.58636e-315
0
7 Pulser~
4 158 73 0 11 12
0 21 167 124 168 0 0 10 10 -1
7 1
0
0 0 4144 0
0
3 V11
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4153 0 0
2
5.89911e-315 5.58669e-315
0
7 74LS126
116 558 241 0 12 25
0 9 97 9 96 9 95 9 94 61
83 82 81
0
0 0 4848 0
7 74LS126
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
8251 0 0
2
5.89911e-315 5.58701e-315
0
7 74LS193
137 393 227 0 14 29
0 124 10 11 130 61 83 82 81 169
170 97 96 95 94
0
0 0 4336 0
7 74LS193
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
8341 0 0
2
5.89911e-315 5.58734e-315
0
7 74LS173
129 598 354 0 14 29
0 2 12 12 124 61 83 82 81 2
2 101 100 99 98
0
0 0 4336 782
7 74LS173
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6192 0 0
2
5.89911e-315 5.58766e-315
0
7 74LS173
129 1253 188 0 14 29
0 2 4 4 124 61 83 82 81 2
2 119 118 117 116
0
0 0 4336 0
7 74LS173
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3842 0 0
2
5.89911e-315 5.58798e-315
0
7 74LS126
116 1103 309 0 12 25
0 5 119 5 118 5 117 5 116 61
83 82 81
0
0 0 4336 512
7 74LS126
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
6185 0 0
2
5.89911e-315 5.58831e-315
0
7 74LS126
116 1105 512 0 12 25
0 2 123 2 122 2 121 2 120 61
83 82 81
0
0 0 4336 512
7 74LS126
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
3914 0 0
2
5.89911e-315 5.58863e-315
0
7 74LS181
132 1249 494 0 22 45
0 6 7 7 6 119 118 117 116 72
73 71 70 7 6 171 172 173 174 123
122 121 120
0
0 0 12528 512
7 74LS181
-24 -69 25 -61
2 U7
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 254
65 0 0 512 1 0 0 0
1 U
367 0 0
2
5.89911e-315 5.58895e-315
0
7 74LS173
129 1272 713 0 14 29
0 2 19 19 124 63 64 65 66 2
2 18 17 16 76
0
0 0 4336 0
7 74LS173
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4366 0 0
2
5.89911e-315 5.58928e-315
0
7 Ground~
168 534 322 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7433 0 0
2
5.89911e-315 5.5896e-315
0
7 Ground~
168 1305 169 0 1 3
0 2
0
0 0 53360 782
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8588 0 0
2
5.89911e-315 5.58993e-315
0
7 Ground~
168 1284 605 0 1 3
0 2
0
0 0 53360 692
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6897 0 0
2
5.89911e-315 5.59025e-315
0
7 74LS157
122 591 517 0 14 29
0 136 98 102 99 103 100 104 101 105
2 106 107 108 109
0
0 0 4336 270
7 74LS157
-24 -60 25 -52
3 U10
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3458 0 0
2
5.89911e-315 5.59057e-315
0
7 Ground~
168 521 503 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5508 0 0
2
5.89911e-315 5.5909e-315
0
6 1K RAM
79 658 666 0 20 41
0 93 93 93 93 93 93 109 108 107
106 88 87 86 85 61 83 82 81 13
20
0
0 0 4336 0
5 RAM1K
-17 -19 18 -11
3 U11
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 1 0 0 0
1 U
3981 0 0
2
5.89911e-315 5.59122e-315
0
7 74LS157
122 708 785 0 14 29
0 135 81 112 82 113 83 114 61 115
2 89 90 111 110
0
0 0 4336 602
7 74LS157
-24 -60 25 -52
3 U12
53 0 74 8
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
4581 0 0
2
5.89911e-315 5.59154e-315
0
7 Ground~
168 626 794 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3346 0 0
2
5.89911e-315 5.59187e-315
0
7 74LS173
129 471 1191 0 14 29
0 2 15 15 124 88 87 86 85 2
2 48 49 50 47
0
0 0 4336 0
7 74LS173
-24 -51 25 -43
3 U13
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
8843 0 0
2
5.89911e-315 5.59219e-315
0
7 Ground~
168 526 1163 0 1 3
0 2
0
0 0 53360 782
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
566 0 0
2
5.89911e-315 5.59252e-315
0
7 Ground~
168 627 1036 0 1 3
0 2
0
0 0 53360 692
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3750 0 0
2
5.89911e-315 5.59284e-315
0
7 74LS173
129 675 1077 0 14 29
0 2 15 15 124 61 83 82 81 14
14 61 83 82 81
0
0 0 4336 0
7 74LS173
-24 -51 25 -43
3 U14
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
9887 0 0
2
5.89911e-315 5.59316e-315
0
14 Logic Display~
6 1420 878 0 1 2
10 132
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
351 0 0
2
5.89911e-315 5.59349e-315
0
14 Logic Display~
6 1443 878 0 1 2
10 131
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7542 0 0
2
5.89911e-315 5.59381e-315
0
14 Logic Display~
6 1397 878 0 1 2
10 133
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9283 0 0
2
5.89911e-315 5.59413e-315
0
14 Logic Display~
6 1374 878 0 1 2
10 134
0
0 0 53360 512
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3600 0 0
2
5.89911e-315 5.59446e-315
0
7 Ground~
168 1293 838 0 1 3
0 2
0
0 0 53360 692
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8274 0 0
2
5.89911e-315 5.59478e-315
0
7 74LS173
129 1255 897 0 14 29
0 2 84 84 124 61 83 82 81 2
2 134 133 132 131
0
0 0 4336 0
7 74LS173
-24 -51 25 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3329 0 0
2
5.89911e-315 5.59511e-315
0
691
1 0 16 0 0 4096 0 37 0 0 215 2
1445 661
1443 661
1 0 17 0 0 4096 0 38 0 0 214 2
1436 639
1436 641
1 0 124 0 0 4096 3 39 0 0 151 2
1435 618
1435 617
1 0 18 0 0 4096 0 40 0 0 213 2
1435 602
1435 601
1 0 19 0 0 4096 0 41 0 0 6 2
1530 519
1530 517
0 0 19 0 0 41088 0 0 0 655 87 12
1217 650
1184 650
1184 581
1464 581
1464 517
1769 517
1769 539
2220 539
2220 570
2874 570
2874 2660
1967 2660
2 0 8 0 0 8192 0 42 0 0 547 3
2357 2200
2357 2202
2464 2202
0 0 20 0 0 4096 0 0 0 144 281 2
143 693
143 713
2 0 11 0 0 16384 0 43 0 0 0 5
2539 2693
2539 2692
2546 2692
2546 2903
2004 2903
1 0 21 0 0 8320 0 364 0 0 156 3
134 64
134 67
110 67
0 0 124 0 0 4096 3 0 0 12 554 3
316 23
787 23
787 67
0 0 124 0 0 0 3 0 0 148 149 2
316 67
316 23
0 0 124 0 0 0 3 0 0 152 553 2
278 242
278 357
0 1 22 0 0 4224 0 0 42 83 0 3
2092 2202
2321 2202
2321 2200
0 0 4 0 0 12288 0 0 0 99 546 8
1692 2642
1750 2642
1750 3040
2535 3040
2535 3056
2739 3056
2739 3050
2761 3050
0 0 5 0 0 8192 0 0 0 82 278 7
2133 2664
2133 2994
2635 2994
2635 3027
2670 3027
2670 3013
2732 3013
0 0 7 0 0 8192 0 0 0 19 275 3
2496 2635
2496 2556
2641 2556
0 0 7 0 0 0 0 0 0 19 162 3
2514 2635
2514 2652
2582 2652
0 0 7 0 0 4096 0 0 0 80 549 2
2240 2635
2551 2635
0 0 14 0 0 4096 0 0 0 91 21 3
1837 2667
1026 2667
1026 2465
0 0 14 0 0 0 0 0 0 280 0 4
226 2428
580 2428
580 2465
1038 2465
0 0 11 0 0 4096 0 0 0 23 545 6
1115 2903
79 2903
79 2764
93 2764
93 2471
86 2471
0 0 11 0 0 0 0 0 0 9 0 2
2007 2903
1110 2903
0 1 23 0 0 4096 0 0 43 39 0 3
2482 2692
2503 2692
2503 2693
0 0 11 0 0 0 0 0 0 545 172 5
86 735
86 357
96 357
96 218
349 218
0 0 6 0 0 4096 0 0 0 77 276 2
2337 2484
2671 2484
0 0 6 0 0 0 0 0 0 77 550 2
2337 2422
2611 2422
0 0 6 0 0 0 0 0 0 77 548 2
2337 2403
2522 2403
0 0 6 0 0 4096 0 0 0 165 548 2
1578 689
2522 689
0 0 13 0 0 4096 0 0 0 31 269 2
543 2268
169 2268
0 0 13 0 0 4096 0 0 0 111 0 4
1492 2376
618 2376
618 2268
540 2268
0 0 15 0 0 4096 0 0 0 119 279 4
1356 2346
642 2346
642 2238
223 2238
0 0 10 0 0 12288 0 0 0 122 544 4
1260 2325
682 2325
682 2211
57 2211
0 0 12 0 0 8192 0 0 0 35 270 3
740 2305
740 2179
114 2179
0 0 12 0 0 0 0 0 0 124 0 2
1142 2305
737 2305
0 0 9 0 0 4096 0 0 0 134 271 2
1100 2090
28 2090
2 0 24 0 0 12288 0 85 0 0 53 4
1770 2344
1770 2339
1733 2339
1733 1861
0 2 25 0 0 4224 0 0 83 110 0 4
1602 2243
1602 2468
1683 2468
1683 2517
0 1 23 0 0 8192 0 0 57 40 0 5
2434 2580
2482 2580
2482 2694
2489 2694
2489 2704
0 1 23 0 0 4224 0 0 61 94 0 5
1919 2434
2434 2434
2434 2637
2431 2637
2431 2677
0 0 26 0 0 4096 0 0 0 97 98 3
1899 2340
1899 2282
1881 2282
0 1 27 0 0 4096 0 0 76 51 0 4
2107 1949
2107 2128
2101 2128
2101 2138
2 0 28 0 0 4096 0 79 0 0 54 2
2054 2456
2054 1836
1 0 29 0 0 4096 0 81 0 0 52 2
1917 2371
1917 1905
1 0 27 0 0 0 0 45 0 0 51 2
1039 1949
1039 1949
1 0 29 0 0 0 0 46 0 0 52 2
1037 1905
1037 1905
1 0 24 0 0 0 0 47 0 0 53 2
1036 1862
1036 1861
1 0 28 0 0 0 0 48 0 0 54 2
1036 1837
1036 1836
1 0 30 0 0 4096 0 49 0 0 55 2
1034 1806
1034 1805
1 0 31 0 0 4096 0 50 0 0 56 2
1024 1776
1024 1775
2 0 27 0 0 4224 0 51 0 0 0 2
1012 1949
2369 1949
2 0 29 0 0 4224 0 52 0 0 0 2
1013 1905
2364 1905
2 0 24 0 0 4224 0 53 0 0 0 2
1023 1861
2383 1861
2 0 28 0 0 4224 0 54 0 0 0 2
1022 1836
2378 1836
2 0 30 0 0 4224 0 55 0 0 0 2
983 1805
2376 1805
2 0 31 0 0 4224 0 56 0 0 0 2
979 1775
2371 1775
17 1 32 0 0 4224 0 96 51 0 0 4
856 1878
927 1878
927 1949
976 1949
18 1 33 0 0 4224 0 96 52 0 0 5
856 1869
945 1869
945 1903
977 1903
977 1905
19 1 34 0 0 4224 0 96 53 0 0 3
856 1860
987 1860
987 1861
20 1 35 0 0 4224 0 96 54 0 0 4
856 1851
958 1851
958 1836
986 1836
21 1 36 0 0 4224 0 96 55 0 0 5
856 1842
917 1842
917 1804
947 1804
947 1805
22 1 37 0 0 8320 0 96 56 0 0 4
856 1833
891 1833
891 1775
943 1775
1 0 38 0 0 4096 0 1 0 0 64 2
702 1510
702 1509
1 0 38 0 0 4224 0 334 0 0 0 2
810 1509
699 1509
1 0 7 0 0 0 0 58 0 0 78 2
2299 2674
2299 2674
1 0 6 0 0 0 0 60 0 0 76 2
2372 2672
2370 2672
1 0 6 0 0 0 0 62 0 0 77 2
2338 2674
2337 2674
1 0 19 0 0 0 0 67 0 0 87 2
1968 2684
1967 2684
1 0 14 0 0 0 0 68 0 0 91 2
1838 2682
1837 2682
1 0 13 0 0 0 0 70 0 0 111 2
1494 2692
1492 2692
1 0 15 0 0 0 0 71 0 0 74 2
1358 2708
1356 2708
1 0 10 0 0 0 0 72 0 0 122 3
1259 2562
1260 2562
1260 2732
1 0 12 0 0 0 0 73 0 0 124 3
1163 2494
1163 2722
1141 2722
0 0 15 0 0 0 0 0 0 119 0 2
1356 2397
1356 2716
0 1 6 0 0 0 0 0 59 76 0 4
2370 2606
2396 2606
2396 2677
2398 2677
0 0 6 0 0 0 0 0 0 77 0 3
2337 2601
2370 2601
2370 2677
0 0 6 0 0 0 0 0 0 104 0 3
1779 2400
2337 2400
2337 2680
0 0 7 0 0 0 0 0 0 79 0 3
2269 2606
2299 2606
2299 2679
0 1 7 0 0 0 0 0 63 80 0 3
2240 2603
2269 2603
2269 2677
0 1 7 0 0 4096 0 0 64 103 0 4
1714 2420
2240 2420
2240 2677
2239 2677
0 1 22 0 0 0 0 0 65 83 0 6
2152 2490
2204 2490
2204 2653
2159 2653
2159 2681
2158 2681
3 1 5 0 0 0 0 75 66 0 0 5
2143 2573
2143 2664
2071 2664
2071 2686
2072 2686
3 1 22 0 0 0 0 76 75 0 0 6
2092 2183
2092 2286
2154 2286
2154 2483
2152 2483
2152 2527
0 2 39 0 0 4224 0 0 75 88 0 3
2064 2510
2134 2510
2134 2527
2 0 26 0 0 0 0 76 0 0 86 3
2083 2138
2084 2138
2084 2098
0 0 26 0 0 4096 0 0 0 513 0 2
2084 1684
2084 2103
2 0 19 0 0 128 0 77 0 0 0 4
2064 2571
2064 2623
1967 2623
1967 2689
1 3 39 0 0 0 0 77 79 0 0 3
2064 2535
2064 2501
2063 2501
1 3 40 0 0 8320 0 78 80 0 0 3
1924 2528
1924 2527
1926 2527
0 1 26 0 0 4096 0 0 79 513 0 5
2030 1684
2030 2307
2087 2307
2087 2456
2072 2456
0 0 14 0 0 0 0 0 0 92 0 2
1837 2603
1837 2687
2 0 14 0 0 0 0 78 0 0 0 3
1924 2564
1924 2603
1826 2603
0 0 41 0 0 4096 0 0 0 0 96 2
1949 2143
1949 2140
3 2 23 0 0 0 0 81 80 0 0 4
1908 2416
1919 2416
1919 2481
1917 2481
0 1 41 0 0 4096 0 0 80 96 0 3
1946 2140
1946 2481
1935 2481
0 0 41 0 0 4224 0 0 0 129 0 2
1151 2140
2010 2140
0 2 26 0 0 0 0 0 81 0 0 2
1899 2334
1899 2371
0 0 26 0 0 0 0 0 0 513 0 4
1853 1684
1853 2087
1881 2087
1881 2339
2 1 4 0 0 0 0 82 69 0 0 3
1692 2599
1692 2678
1690 2678
1 3 42 0 0 0 0 82 83 0 0 2
1692 2563
1692 2563
3 1 43 0 0 8320 0 84 83 0 0 4
1724 2486
1724 2506
1701 2506
1701 2517
2 0 7 0 0 0 0 84 0 0 103 2
1715 2440
1714 2440
3 0 7 0 0 0 0 86 0 0 0 4
1672 2367
1672 2420
1714 2420
1714 2444
3 1 6 0 0 0 0 85 84 0 0 4
1779 2389
1779 2416
1733 2416
1733 2440
1 0 26 0 0 0 0 85 0 0 106 2
1788 2344
1790 2344
0 0 26 0 0 0 0 0 0 107 0 7
1699 2237
1836 2237
1836 2307
1771 2307
1771 2333
1790 2333
1790 2349
0 1 26 0 0 0 0 0 86 513 0 4
1699 1684
1699 2283
1681 2283
1681 2322
2 0 30 0 0 0 0 86 0 0 109 2
1663 2322
1664 2322
0 0 30 0 0 0 0 0 0 55 0 2
1664 1805
1664 2330
0 0 25 0 0 0 0 0 0 115 0 2
1500 2243
1640 2243
2 0 13 0 0 0 0 87 0 0 0 2
1492 2337
1492 2696
1 3 44 0 0 4224 0 87 88 0 0 3
1492 2301
1492 2303
1491 2303
0 0 10 0 0 0 0 0 0 118 114 3
1443 2104
1469 2104
1469 2117
0 2 10 0 0 0 0 0 88 0 0 4
1469 2111
1469 2224
1482 2224
1482 2257
3 1 25 0 0 0 0 89 88 0 0 4
1495 2220
1495 2235
1500 2235
1500 2257
0 1 45 0 0 4096 0 0 89 527 0 3
1519 1712
1519 2175
1504 2175
0 2 31 0 0 0 0 0 89 56 0 3
1487 1775
1487 2175
1486 2175
0 0 10 0 0 0 0 0 0 122 0 2
1260 2104
1466 2104
2 0 15 0 0 0 0 90 0 0 0 2
1356 2261
1356 2401
1 0 10 0 0 0 0 90 0 0 121 2
1356 2225
1356 2225
0 0 10 0 0 0 0 0 0 122 0 3
1260 2146
1356 2146
1356 2229
0 0 10 0 0 4096 0 0 0 528 0 2
1260 1654
1260 2736
0 0 10 0 0 0 0 0 0 528 528 2
1188 1654
1241 1654
2 0 12 0 0 0 0 91 0 0 0 4
1142 2282
1142 2716
1141 2716
1141 2726
1 0 46 0 0 0 0 91 0 0 126 2
1142 2246
1142 2246
3 0 46 0 0 4224 0 92 0 0 0 2
1142 2207
1142 2250
0 1 9 0 0 0 0 0 74 134 0 3
1100 2164
1100 2733
1099 2733
0 2 9 0 0 0 0 0 92 134 0 3
1100 2036
1133 2036
1133 2161
1 3 41 0 0 0 0 92 93 0 0 4
1151 2161
1151 2140
1157 2140
1157 2131
2 0 26 0 0 0 0 93 0 0 133 2
1148 2086
1149 2086
1 0 31 0 0 0 0 93 0 0 132 2
1166 2086
1164 2086
0 0 31 0 0 0 0 0 0 56 0 2
1164 1775
1164 2091
0 0 26 0 0 0 0 0 0 513 0 2
1149 1684
1149 2091
0 0 9 0 0 0 0 0 0 529 0 2
1100 1627
1100 2172
1 0 2 0 0 4096 0 95 0 0 136 2
588 1921
588 1923
0 0 2 0 0 4096 0 0 0 137 0 2
726 1923
583 1923
1 2 2 0 0 0 0 96 96 0 0 4
780 1923
721 1923
721 1914
780 1914
0 1 47 0 0 4096 0 0 5 143 0 2
570 1860
539 1860
1 0 48 0 0 4096 0 2 0 0 140 4
469 1892
525 1892
525 1887
550 1887
3 0 48 0 0 4096 0 96 0 0 0 2
786 1887
544 1887
4 1 49 0 0 4096 0 96 3 0 0 4
786 1878
508 1878
508 1881
493 1881
5 1 50 0 0 4096 0 96 4 0 0 4
786 1869
540 1869
540 1871
513 1871
6 1 47 0 0 4096 0 96 5 0 0 2
786 1860
539 1860
0 20 20 0 0 16512 0 0 378 0 0 9
143 701
143 662
141 662
141 644
501 644
501 591
708 591
708 639
696 639
0 2 20 0 0 0 0 0 97 144 0 2
395 644
395 850
0 3 4 0 0 0 0 0 368 0 0 4
1620 108
1167 108
1167 179
1215 179
0 0 51 0 0 4224 0 0 0 0 0 2
1632 108
1624 108
0 0 124 0 0 0 3 0 0 0 262 2
316 48
316 67
0 0 124 0 0 0 3 0 0 0 0 2
316 23
316 44
0 0 52 0 0 4224 0 0 0 0 0 2
386 23
386 34
0 4 124 0 0 0 3 0 108 555 0 4
1417 617
1750 617
1750 642
1804 642
0 0 124 0 0 0 3 0 0 0 262 2
278 257
278 200
1 0 124 0 0 0 3 98 0 0 230 2
737 68
737 67
1 0 53 0 0 4224 0 6 0 0 0 4
511 56
524 56
524 65
536 65
0 1 53 0 0 0 0 0 6 0 0 2
516 56
511 56
1 0 21 0 0 0 0 26 0 0 0 2
101 67
114 67
0 1 21 0 0 0 0 0 26 0 0 2
106 67
101 67
2 0 13 0 0 0 0 99 0 0 647 2
443 706
443 673
1 1 54 0 0 8320 0 7 99 0 0 3
473 722
477 722
477 706
0 0 55 0 0 4096 0 0 0 0 0 3
1730 550
1730 634
1811 634
1 0 56 0 0 4096 0 17 0 0 0 2
1631 108
1628 108
0 2 7 0 0 4224 0 0 371 0 0 7
2582 2846
2582 456
1877 456
1877 453
1852 453
1852 458
1281 458
0 0 57 0 0 4224 0 0 0 0 0 3
1887 452
1882 452
1882 456
0 1 6 0 0 0 0 0 371 0 0 4
1861 417
1856 417
1856 449
1281 449
0 1 6 0 0 0 0 0 106 0 0 3
1585 689
1568 689
1568 721
0 0 45 0 0 0 0 0 0 527 527 2
1269 1712
1273 1712
0 2 10 0 0 0 0 0 366 282 0 4
69 239
69 208
361 208
361 209
0 1 58 0 0 4224 0 0 18 0 0 2
223 1286
223 1295
0 0 14 0 0 0 0 0 0 0 280 5
196 1106
196 1091
180 1091
180 1204
196 1204
0 0 13 0 0 0 0 0 0 0 263 3
177 748
168 748
168 735
0 0 55 0 0 12416 0 0 0 160 0 5
1730 564
1642 564
1642 589
1500 589
1500 584
3 0 11 0 0 0 0 366 0 0 0 2
355 218
345 218
3 1 59 0 0 8320 0 104 102 0 0 4
388 801
388 802
420 802
420 799
2 2 60 0 0 4224 0 103 104 0 0 2
324 810
343 810
0 1 61 0 0 16384 0 0 104 560 0 7
1066 494
1066 472
736 472
736 400
330 400
330 792
343 792
0 0 9 0 0 0 0 0 0 529 0 2
1014 1627
1014 1639
0 0 10 0 0 0 0 0 0 528 0 2
994 1654
994 1674
0 0 49 0 0 0 0 0 0 536 141 4
528 1662
528 1787
745 1787
745 1878
1 8 62 0 0 12416 0 8 108 0 0 5
1803 1001
1803 1002
1790 1002
1790 678
1804 678
5 1 63 0 0 4224 0 372 9 0 0 6
1240 722
1157 722
1157 642
1076 642
1076 671
1090 671
6 1 64 0 0 12416 0 372 10 0 0 6
1240 731
1164 731
1164 721
1082 721
1082 706
1086 706
7 1 65 0 0 12416 0 372 11 0 0 5
1240 740
1179 740
1179 761
1086 761
1086 745
8 1 66 0 0 12416 0 372 12 0 0 5
1240 749
1198 749
1198 791
1084 791
1084 782
1 5 67 0 0 8320 0 14 108 0 0 4
1823 866
1762 866
1762 651
1804 651
1 6 68 0 0 8320 0 15 108 0 0 4
1823 900
1773 900
1773 660
1804 660
1 7 69 0 0 8320 0 13 108 0 0 4
1823 942
1783 942
1783 669
1804 669
0 0 8 0 0 8192 0 0 0 0 547 4
1656 814
1656 847
2104 847
2104 814
0 0 4 0 0 0 0 0 0 546 146 4
1903 108
1903 40
1567 40
1567 108
0 0 6 0 0 0 0 0 0 272 548 4
1863 543
1863 564
2132 564
2132 476
0 0 6 0 0 0 0 0 0 272 272 2
1877 543
1880 543
0 0 7 0 0 0 0 0 0 267 549 6
1882 499
1882 523
2043 523
2043 495
2088 495
2088 467
0 0 7 0 0 0 0 0 0 552 275 4
1648 401
1648 187
2021 187
2021 401
0 0 6 0 0 0 0 0 0 551 276 4
1672 381
1672 288
1925 288
1925 381
0 0 6 0 0 0 0 0 0 551 551 2
1692 381
1685 381
0 0 2 0 0 8192 0 0 0 0 277 4
1896 362
1896 312
1711 312
1711 362
0 0 5 0 0 0 0 0 0 278 673 4
1901 270
1901 215
1694 215
1694 270
0 0 15 0 0 0 0 0 0 279 507 4
223 1352
254 1352
254 1276
223 1276
0 0 12 0 0 0 0 0 0 270 264 3
114 386
151 386
151 304
0 0 10 0 0 0 0 0 0 544 167 5
57 338
74 338
74 258
88 258
88 208
0 0 9 0 0 0 0 0 0 271 542 5
28 325
7 325
7 81
84 81
84 108
0 0 48 0 0 4096 0 0 0 537 140 4
537 1521
537 1807
736 1807
736 1887
2 0 55 0 0 0 0 108 0 0 160 3
1798 624
1782 624
1782 634
1 0 2 0 0 0 0 108 0 0 223 4
1804 615
1787 615
1787 590
1895 590
10 0 2 0 0 0 0 108 0 0 223 3
1874 624
1895 624
1895 614
12 0 70 0 0 0 0 371 0 0 210 2
1287 548
1287 548
11 0 71 0 0 0 0 371 0 0 209 2
1287 539
1287 539
14 9 72 0 0 8320 0 106 371 0 0 4
1496 785
1360 785
1360 521
1287 521
13 10 73 0 0 12416 0 106 371 0 0 5
1514 785
1514 822
1348 822
1348 530
1287 530
12 0 71 0 0 12416 0 106 0 0 0 5
1532 785
1532 839
1335 839
1335 539
1284 539
11 0 70 0 0 12416 0 106 0 0 0 5
1550 785
1550 829
1324 829
1324 548
1283 548
0 0 74 0 0 4224 0 0 0 0 0 2
1597 689
1589 689
10 0 75 0 0 8320 0 106 0 0 0 3
1487 715
1453 715
1453 762
11 9 18 0 0 8320 0 372 106 0 0 5
1304 722
1388 722
1388 601
1496 601
1496 721
12 7 17 0 0 4224 0 372 106 0 0 5
1304 731
1431 731
1431 641
1514 641
1514 721
13 5 16 0 0 4224 0 372 106 0 0 5
1304 740
1443 740
1443 661
1532 661
1532 721
14 3 76 0 0 4224 0 372 106 0 0 5
1304 749
1456 749
1456 690
1550 690
1550 721
6 0 77 0 0 4096 0 106 0 0 220 4
1523 721
1523 694
1532 694
1532 679
4 0 78 0 0 4096 0 106 0 0 221 4
1541 721
1541 694
1550 694
1550 679
11 8 79 0 0 12416 0 108 106 0 0 7
1868 651
1934 651
1934 701
1679 701
1679 608
1505 608
1505 721
12 0 77 0 0 12416 0 108 0 0 0 7
1868 660
1903 660
1903 721
1660 721
1660 629
1532 629
1532 683
13 0 78 0 0 12416 0 108 0 0 0 7
1868 669
1916 669
1916 743
1643 743
1643 639
1550 639
1550 684
14 2 80 0 0 12416 0 108 106 0 0 7
1868 678
1890 678
1890 759
1629 759
1629 654
1559 654
1559 721
1 9 2 0 0 0 0 107 108 0 0 3
1895 578
1895 615
1874 615
0 0 81 0 0 4096 0 0 0 538 254 2
443 161
484 161
0 0 82 0 0 4096 0 0 0 539 255 2
443 154
483 154
0 0 83 0 0 4096 0 0 0 540 256 2
442 146
483 146
0 0 61 0 0 0 0 0 0 541 257 2
442 138
482 138
0 3 84 0 0 4224 0 0 390 0 0 4
1660 814
1189 814
1189 888
1217 888
1 0 56 0 0 4224 0 17 0 0 0 2
1631 108
1626 108
0 0 124 0 0 0 3 0 0 0 554 3
596 65
596 67
737 67
0 0 85 0 0 4096 0 0 0 238 258 2
867 441
867 420
0 0 86 0 0 4096 0 0 0 239 259 2
836 437
836 418
0 0 85 0 0 4096 0 0 0 688 238 2
867 792
867 770
0 0 86 0 0 0 0 0 0 689 239 2
836 793
836 774
0 0 87 0 0 4096 0 0 0 690 240 2
804 793
804 772
0 0 88 0 0 4096 0 0 0 691 241 2
772 790
772 774
0 2 124 0 0 0 3 0 229 412 0 4
278 1302
357 1302
357 1470
724 1470
0 0 85 0 0 4096 0 0 0 0 0 2
867 778
867 433
0 0 86 0 0 4096 0 0 0 0 0 2
836 779
836 428
0 0 87 0 0 4096 0 0 0 0 260 2
804 780
804 423
0 0 88 0 0 4096 0 0 0 0 0 2
772 780
772 428
0 15 61 0 0 0 0 0 378 0 0 3
697 715
697 684
690 684
0 16 83 0 0 0 0 0 378 0 0 3
702 718
702 693
690 693
0 17 82 0 0 0 0 0 378 0 0 3
707 716
707 702
690 702
0 18 81 0 0 0 0 0 378 0 0 3
725 715
725 711
690 711
11 0 89 0 0 4224 0 379 0 0 0 2
725 752
725 719
0 0 61 0 0 0 0 0 0 249 596 2
790 684
779 684
12 0 90 0 0 4224 0 379 0 0 0 2
707 752
707 720
0 0 61 0 0 0 0 0 0 0 687 2
787 684
924 684
0 0 83 0 0 4096 0 0 0 0 686 2
790 693
954 693
0 0 82 0 0 4096 0 0 0 0 684 2
788 702
984 702
0 0 81 0 0 4096 0 0 0 0 685 2
791 711
1013 711
0 0 124 0 0 0 3 0 0 0 613 2
278 351
278 297
0 0 81 0 0 4096 0 0 0 0 685 2
460 161
1013 161
0 0 82 0 0 4096 0 0 0 0 684 2
461 154
984 154
0 0 83 0 0 4096 0 0 0 0 686 2
463 146
954 146
0 0 61 0 0 4096 0 0 0 0 687 2
465 138
924 138
0 0 85 0 0 0 0 0 0 0 0 2
867 429
867 130
0 0 86 0 0 0 0 0 0 0 0 2
836 424
836 131
0 0 87 0 0 0 0 0 0 0 0 2
804 429
804 132
0 0 88 0 0 0 0 0 0 241 0 2
772 431
772 132
1 0 124 0 0 0 3 366 0 0 0 4
361 200
278 200
278 67
361 67
1 0 13 0 0 0 0 322 0 0 0 3
174 673
168 673
168 739
0 0 12 0 0 0 0 0 0 266 0 4
151 304
112 304
112 303
68 303
2 1 12 0 0 0 0 367 320 0 0 3
578 318
578 304
178 304
0 1 12 0 0 0 0 0 320 0 0 2
148 304
178 304
0 0 7 0 0 0 0 0 0 0 273 4
1892 499
1873 499
1873 467
1847 467
1 0 91 0 0 4224 0 19 0 0 0 2
196 1115
196 1110
0 1 13 0 0 16512 0 0 349 263 0 5
168 731
221 731
221 827
169 827
169 2455
0 1 12 0 0 4224 0 0 348 0 0 2
114 365
114 2585
0 1 9 0 0 4224 0 0 345 0 0 2
28 315
28 2768
0 4 6 0 0 0 0 0 371 0 0 4
1890 543
1856 543
1856 476
1281 476
0 3 7 0 0 0 0 0 371 0 0 2
1854 467
1281 467
1 0 92 0 0 4224 0 16 0 0 0 2
1875 417
1865 417
0 1 7 0 0 0 0 0 339 0 0 3
1892 401
2641 401
2641 2785
0 1 6 0 0 8320 0 0 338 0 0 3
1894 381
2671 381
2671 2857
1 1 2 0 0 16512 0 44 370 0 0 7
1750 366
1750 361
1722 361
1722 362
1166 362
1166 485
1137 485
0 1 5 0 0 8320 0 0 336 0 0 3
1896 270
2732 270
2732 3024
0 1 15 0 0 4224 0 0 351 0 0 2
223 1347
223 2339
0 1 14 0 0 4224 0 0 350 0 0 4
196 1197
196 2381
226 2381
226 2458
1 0 20 0 0 0 0 20 0 0 0 2
143 755
143 705
0 0 10 0 0 0 0 0 0 0 0 4
45 240
45 239
69 239
69 217
1 1 93 0 0 4224 0 22 378 0 0 2
626 583
626 630
2 1 93 0 0 0 0 378 378 0 0 2
626 639
626 630
3 2 93 0 0 0 0 378 378 0 0 2
626 648
626 639
4 3 93 0 0 0 0 378 378 0 0 2
626 657
626 648
5 4 93 0 0 0 0 378 378 0 0 2
626 666
626 657
6 5 93 0 0 0 0 378 378 0 0 2
626 675
626 666
1 0 81 0 0 0 0 109 0 0 685 2
1013 1350
1013 1350
1 0 82 0 0 0 0 110 0 0 684 2
984 1350
984 1350
1 0 83 0 0 0 0 111 0 0 686 2
954 1350
954 1350
1 0 61 0 0 0 0 112 0 0 687 2
924 1350
924 1350
1 0 85 0 0 0 0 113 0 0 688 2
867 1350
867 1350
1 0 86 0 0 0 0 114 0 0 689 2
836 1350
836 1350
1 0 87 0 0 0 0 115 0 0 690 2
804 1349
804 1349
1 0 88 0 0 0 0 116 0 0 691 2
772 1349
772 1349
1 0 88 0 0 0 0 117 0 0 691 2
772 980
772 980
1 0 87 0 0 0 0 118 0 0 690 2
804 980
804 980
1 0 86 0 0 0 0 119 0 0 689 2
836 980
836 980
1 0 85 0 0 0 0 120 0 0 688 2
867 980
867 980
1 0 61 0 0 0 0 121 0 0 687 2
924 980
924 980
1 0 83 0 0 0 0 122 0 0 686 2
954 980
954 980
1 0 82 0 0 0 0 123 0 0 684 2
984 980
984 980
1 0 81 0 0 0 0 124 0 0 685 2
1013 979
1013 979
1 0 88 0 0 0 0 125 0 0 241 2
772 604
772 604
1 0 87 0 0 0 0 126 0 0 240 2
804 604
804 604
1 0 86 0 0 0 0 127 0 0 239 2
836 603
836 603
1 0 85 0 0 0 0 128 0 0 238 2
867 603
867 603
1 0 61 0 0 0 0 129 0 0 687 2
924 604
924 604
1 0 83 0 0 0 0 130 0 0 686 2
954 604
954 604
1 0 82 0 0 0 0 131 0 0 684 2
984 604
984 604
1 0 81 0 0 0 0 132 0 0 685 2
1013 604
1013 604
1 0 81 0 0 0 0 133 0 0 605 2
597 277
597 277
1 0 82 0 0 0 0 134 0 0 606 2
597 259
597 259
1 0 83 0 0 0 0 135 0 0 607 2
597 241
597 241
1 0 61 0 0 0 0 136 0 0 608 2
597 223
597 223
1 0 94 0 0 0 0 137 0 0 678 2
473 277
473 277
1 0 95 0 0 0 0 138 0 0 679 2
473 259
473 259
1 0 96 0 0 0 0 139 0 0 680 2
473 241
473 241
1 0 97 0 0 0 0 140 0 0 677 2
473 223
473 223
1 0 81 0 0 0 0 141 0 0 538 2
335 263
335 263
1 0 82 0 0 0 0 142 0 0 539 3
321 253
321 254
327 254
1 0 83 0 0 0 0 143 0 0 540 2
304 245
318 245
1 0 61 0 0 0 0 144 0 0 541 2
290 236
309 236
1 0 81 0 0 0 0 145 0 0 601 3
736 349
742 349
742 350
1 0 82 0 0 0 0 146 0 0 602 3
714 331
719 331
719 332
1 0 83 0 0 0 0 147 0 0 603 2
687 312
695 312
1 0 61 0 0 0 0 148 0 0 604 3
663 296
672 296
672 297
1 0 98 0 0 0 0 149 0 0 609 2
617 432
617 432
1 0 99 0 0 0 0 150 0 0 610 2
599 423
599 423
1 0 100 0 0 4096 0 151 0 0 611 2
581 413
581 414
1 0 101 0 0 0 0 152 0 0 612 2
563 406
563 406
1 0 102 0 0 0 0 153 0 0 649 2
462 510
462 510
1 0 103 0 0 0 0 154 0 0 650 2
434 510
434 510
1 0 104 0 0 0 0 155 0 0 651 2
405 510
405 510
1 0 105 0 0 0 0 156 0 0 652 2
374 510
374 510
1 0 106 0 0 0 0 157 0 0 643 2
608 621
608 621
1 0 107 0 0 0 0 158 0 0 644 2
590 621
590 621
1 0 108 0 0 4096 0 159 0 0 645 2
572 621
572 622
1 0 109 0 0 0 0 160 0 0 646 2
554 621
554 621
1 0 81 0 0 0 0 161 0 0 593 2
759 711
759 711
1 0 82 0 0 0 0 162 0 0 594 2
759 702
759 702
1 0 83 0 0 0 0 163 0 0 595 2
759 693
759 693
1 0 61 0 0 0 0 164 0 0 596 2
759 684
759 684
1 0 85 0 0 0 0 165 0 0 597 2
759 675
759 675
1 0 86 0 0 0 0 166 0 0 598 2
759 666
759 666
1 0 87 0 0 0 0 167 0 0 599 2
759 657
759 657
1 0 88 0 0 0 0 168 0 0 600 2
759 648
759 648
1 2 81 0 0 0 0 173 379 0 0 4
734 867
734 813
734 813
734 816
1 4 82 0 0 0 0 174 379 0 0 4
716 867
716 813
716 813
716 816
1 6 83 0 0 0 0 175 379 0 0 4
698 868
698 814
698 814
698 816
1 8 61 0 0 0 0 176 379 0 0 4
680 868
680 813
680 813
680 816
1 11 89 0 0 0 0 169 379 0 0 2
725 756
725 752
1 12 90 0 0 0 0 170 379 0 0 2
707 756
707 752
1 14 110 0 0 4096 0 171 379 0 0 2
671 756
671 752
1 13 111 0 0 4096 0 172 379 0 0 2
689 755
689 752
1 0 112 0 0 0 0 177 0 0 633 2
540 892
540 892
1 0 113 0 0 0 0 178 0 0 634 2
512 892
512 892
1 0 114 0 0 0 0 179 0 0 635 2
484 892
484 892
1 0 115 0 0 0 0 180 0 0 636 2
452 892
452 892
1 0 81 0 0 0 0 181 0 0 585 2
719 1161
719 1161
1 0 82 0 0 0 0 182 0 0 586 2
698 1152
698 1152
1 0 83 0 0 0 0 183 0 0 587 2
679 1143
679 1143
1 0 61 0 0 0 0 184 0 0 588 2
660 1134
660 1134
1 0 85 0 0 0 0 185 0 0 589 2
485 1277
485 1277
1 0 86 0 0 0 0 186 0 0 590 2
471 1267
471 1267
1 0 87 0 0 0 0 187 0 0 591 2
460 1258
460 1258
1 0 88 0 0 0 0 188 0 0 592 2
449 1248
449 1248
1 0 47 0 0 0 0 189 0 0 534 2
510 1343
510 1343
1 0 50 0 0 0 0 190 0 0 535 2
519 1322
519 1322
1 0 49 0 0 0 0 191 0 0 536 2
528 1301
528 1301
1 0 48 0 0 0 0 192 0 0 537 2
538 1285
537 1285
1 0 81 0 0 0 0 193 0 0 618 2
742 1113
742 1113
1 0 82 0 0 0 0 194 0 0 619 2
735 1104
735 1104
1 0 83 0 0 0 0 195 0 0 620 2
724 1095
724 1095
1 0 61 0 0 0 0 196 0 0 621 2
711 1086
711 1086
1 0 81 0 0 0 0 197 0 0 557 2
1060 548
1060 548
1 0 82 0 0 0 0 198 0 0 558 2
1060 530
1060 530
1 0 83 0 0 0 0 199 0 0 559 2
1060 512
1060 512
1 0 61 0 0 0 0 200 0 0 560 2
1060 494
1060 494
1 0 81 0 0 0 0 201 0 0 581 2
1060 345
1060 345
1 0 82 0 0 0 0 202 0 0 582 2
1060 327
1060 327
1 0 83 0 0 0 0 203 0 0 583 2
1060 309
1060 309
1 0 61 0 0 0 0 204 0 0 584 2
1060 291
1060 291
1 0 116 0 0 4096 0 205 0 0 669 2
1184 346
1184 345
1 0 117 0 0 0 0 206 0 0 670 2
1184 327
1184 327
1 0 118 0 0 0 0 207 0 0 671 2
1184 309
1184 309
1 0 119 0 0 0 0 208 0 0 672 2
1183 291
1183 291
1 0 120 0 0 0 0 209 0 0 662 2
1160 548
1160 548
1 0 121 0 0 0 0 210 0 0 663 2
1160 530
1160 530
1 0 122 0 0 0 0 211 0 0 664 2
1160 512
1160 512
1 0 123 0 0 0 0 212 0 0 665 2
1160 494
1160 494
1 0 116 0 0 0 0 213 0 0 658 2
1349 413
1349 413
1 0 117 0 0 0 0 214 0 0 659 2
1335 413
1335 413
1 0 118 0 0 0 0 215 0 0 660 2
1321 413
1321 413
1 0 119 0 0 0 0 216 0 0 661 2
1308 413
1308 413
1 0 116 0 0 0 0 217 0 0 669 2
1349 231
1349 231
1 0 117 0 0 0 0 218 0 0 670 2
1335 231
1335 231
1 0 118 0 0 0 0 219 0 0 671 2
1321 231
1321 231
1 0 119 0 0 0 0 220 0 0 672 2
1308 231
1308 231
1 0 81 0 0 0 0 221 0 0 561 2
1114 933
1114 933
1 0 82 0 0 0 0 222 0 0 562 2
1093 924
1093 924
1 0 83 0 0 0 0 223 0 0 563 2
1070 915
1070 915
1 0 61 0 0 0 0 224 0 0 564 2
1050 905
1050 906
1 0 81 0 0 0 0 225 0 0 573 2
1110 224
1110 224
1 0 82 0 0 0 0 226 0 0 574 2
1086 215
1086 215
1 0 83 0 0 0 0 227 0 0 575 2
1061 206
1061 206
1 0 61 0 0 0 0 228 0 0 576 2
1040 197
1040 197
3 0 124 0 0 4096 0 334 0 0 410 3
858 1509
914 1509
914 1470
1 3 124 0 0 4224 0 229 362 0 0 2
758 1470
1176 1470
1 0 124 0 0 0 3 230 0 0 237 2
648 1470
648 1470
4 0 124 0 0 8320 3 381 0 0 0 4
439 1191
278 1191
278 2307
327 2307
1 0 4 0 0 0 0 231 0 0 546 2
2761 3083
2761 3083
1 0 5 0 0 0 0 232 0 0 278 2
2732 2996
2732 2996
1 0 6 0 0 0 0 234 0 0 276 2
2671 2838
2671 2838
1 0 7 0 0 0 0 235 0 0 275 2
2641 2764
2641 2764
1 0 6 0 0 0 0 236 0 0 550 2
2611 2688
2611 2688
1 0 7 0 0 0 0 238 0 0 549 2
2551 2548
2551 2548
1 0 6 0 0 0 0 239 0 0 548 2
2522 2466
2522 2466
1 0 8 0 0 0 0 240 0 0 547 2
2463 2308
2464 2308
1 0 4 0 0 0 0 241 0 0 546 2
2762 2276
2761 2276
1 0 5 0 0 0 0 242 0 0 278 2
2731 2254
2732 2254
1 0 6 0 0 0 0 244 0 0 276 2
2671 2206
2671 2206
1 0 7 0 0 0 0 245 0 0 275 2
2642 2186
2641 2186
1 0 6 0 0 0 0 246 0 0 550 2
2612 2158
2611 2158
1 0 7 0 0 0 0 248 0 0 549 2
2551 2118
2551 2118
1 0 6 0 0 0 0 249 0 0 548 2
2522 2092
2522 2092
1 0 8 0 0 0 0 250 0 0 547 2
2463 2036
2464 2036
1 0 4 0 0 0 0 251 0 0 546 2
2761 1748
2761 1748
1 0 5 0 0 0 0 252 0 0 278 2
2732 1732
2732 1732
1 0 6 0 0 0 0 253 0 0 276 2
2670 1696
2671 1696
1 0 7 0 0 0 0 254 0 0 275 2
2641 1680
2641 1680
1 0 6 0 0 0 0 255 0 0 550 2
2611 1668
2611 1668
1 0 7 0 0 0 0 257 0 0 549 2
2551 1636
2551 1636
1 0 6 0 0 0 0 258 0 0 548 2
2522 1616
2522 1616
1 0 8 0 0 0 0 259 0 0 437 2
2463 1549
2463 1549
1 0 8 0 0 0 0 260 0 0 547 2
2463 1549
2464 1549
1 0 4 0 0 0 0 261 0 0 546 2
2762 1325
2761 1325
1 0 5 0 0 0 0 262 0 0 278 2
2733 1304
2732 1304
1 0 6 0 0 0 0 263 0 0 276 2
2671 1269
2671 1269
1 0 7 0 0 0 0 264 0 0 275 2
2642 1248
2641 1248
1 0 6 0 0 0 0 265 0 0 550 2
2612 1222
2611 1222
1 0 7 0 0 0 0 267 0 0 549 2
2551 1188
2551 1188
1 0 6 0 0 0 0 268 0 0 548 2
2522 1170
2522 1170
1 0 8 0 0 0 0 269 0 0 547 2
2463 1131
2464 1131
1 0 4 0 0 0 0 270 0 0 546 2
2761 562
2761 562
1 0 5 0 0 0 0 271 0 0 278 2
2732 538
2732 538
1 0 6 0 0 0 0 272 0 0 276 2
2671 488
2671 488
1 0 7 0 0 0 0 273 0 0 275 2
2641 468
2641 468
1 0 6 0 0 0 0 274 0 0 550 2
2611 566
2611 566
1 0 7 0 0 0 0 276 0 0 549 2
2551 537
2551 537
1 0 6 0 0 0 0 277 0 0 548 2
2522 523
2522 523
1 0 4 0 0 0 0 278 0 0 546 2
2761 921
2761 921
1 0 5 0 0 0 0 279 0 0 278 2
2732 900
2732 900
1 0 6 0 0 0 0 280 0 0 276 2
2671 865
2671 865
1 0 7 0 0 0 0 281 0 0 275 2
2641 842
2641 842
1 0 6 0 0 0 0 282 0 0 550 2
2611 816
2611 816
1 0 7 0 0 0 0 284 0 0 549 2
2552 773
2551 773
1 0 6 0 0 0 0 285 0 0 548 2
2522 750
2522 750
1 0 9 0 0 0 0 286 0 0 271 2
27 2756
28 2756
1 0 10 0 0 0 0 287 0 0 544 2
57 2698
57 2698
1 0 11 0 0 0 0 288 0 0 545 2
85 2634
86 2634
1 0 12 0 0 0 0 289 0 0 270 2
113 2570
114 2570
1 0 13 0 0 0 0 290 0 0 269 2
169 2442
169 2442
1 0 14 0 0 0 0 291 0 0 280 2
196 2381
196 2381
1 0 15 0 0 0 0 292 0 0 279 2
223 2327
223 2327
1 0 15 0 0 0 0 293 0 0 279 2
224 2062
223 2062
1 0 14 0 0 0 0 294 0 0 280 2
196 2015
196 2015
1 0 13 0 0 0 0 295 0 0 269 2
169 1967
169 1967
1 0 12 0 0 0 0 296 0 0 270 2
113 1850
114 1850
1 0 11 0 0 0 0 297 0 0 545 2
86 1794
86 1794
1 0 10 0 0 0 0 298 0 0 544 2
57 1744
57 1744
1 0 9 0 0 0 0 299 0 0 271 2
28 1704
28 1704
1 0 15 0 0 0 0 300 0 0 279 2
223 1450
223 1450
1 0 14 0 0 0 0 301 0 0 280 2
196 1394
196 1394
1 0 13 0 0 0 0 302 0 0 269 2
169 1348
169 1348
1 0 12 0 0 0 0 303 0 0 270 2
115 1266
114 1266
1 0 11 0 0 0 0 304 0 0 545 2
85 1230
86 1230
1 0 10 0 0 0 0 305 0 0 544 2
57 1184
57 1184
1 0 9 0 0 0 0 306 0 0 271 2
28 1140
28 1140
1 0 15 0 0 0 0 307 0 0 507 2
223 1191
223 1191
1 0 14 0 0 0 0 308 0 0 506 2
196 1026
196 1026
1 0 13 0 0 0 0 309 0 0 269 2
169 924
169 924
1 0 12 0 0 0 0 310 0 0 270 2
114 842
114 842
1 0 11 0 0 0 0 311 0 0 545 2
86 788
86 788
1 0 10 0 0 0 0 312 0 0 544 2
57 749
57 749
1 0 9 0 0 0 0 313 0 0 271 2
28 725
28 725
1 0 12 0 0 0 0 314 0 0 270 2
114 536
114 536
1 0 10 0 0 0 0 315 0 0 544 2
57 448
57 448
1 0 9 0 0 0 0 316 0 0 271 2
28 414
28 414
1 0 9 0 0 0 0 317 0 0 542 4
517 108
516 108
516 109
515 109
1 0 9 0 0 0 0 318 0 0 542 2
179 107
179 108
1 0 10 0 0 0 0 319 0 0 167 2
144 209
144 208
1 0 20 0 0 0 0 321 0 0 144 2
174 644
174 644
1 0 84 0 0 0 0 323 0 0 228 2
1634 813
1634 814
1 0 6 0 0 0 0 325 0 0 272 2
1744 476
1744 476
1 0 7 0 0 0 0 326 0 0 273 2
1707 467
1707 467
1 0 7 0 0 0 0 327 0 0 162 2
1665 458
1665 458
1 0 6 0 0 0 0 328 0 0 164 2
1625 448
1625 449
1 0 7 0 0 0 0 329 0 0 552 2
1625 400
1625 401
1 0 6 0 0 0 0 330 0 0 551 2
1625 380
1625 381
1 0 2 0 0 0 0 331 0 0 277 2
1625 361
1625 362
1 0 5 0 0 0 0 332 0 0 673 2
1622 269
1622 270
1 0 4 0 0 0 0 333 0 0 146 2
1617 108
1617 108
1 0 38 0 0 0 0 334 0 0 0 2
810 1509
806 1509
9 0 14 0 0 0 0 384 0 0 169 5
713 1050
714 1050
714 1026
196 1026
196 1092
2 0 15 0 0 0 0 381 0 0 0 3
433 1173
223 1173
223 1282
1 0 9 0 0 0 0 352 0 0 529 2
911 1627
911 1627
1 0 10 0 0 0 0 353 0 0 528 2
911 1654
911 1654
1 0 26 0 0 0 0 354 0 0 513 2
911 1684
911 1684
1 0 45 0 0 0 0 355 0 0 527 2
911 1712
911 1712
0 1 125 0 0 4096 0 0 25 524 0 2
1168 1528
1069 1528
9 1 26 0 0 20608 0 362 357 0 0 6
1246 1461
1263 1461
1263 1599
798 1599
798 1684
2272 1684
12 2 126 0 0 12416 0 361 362 0 0 6
1477 1503
1521 1503
1521 1373
1118 1373
1118 1461
1182 1461
11 1 10 0 0 0 0 361 362 0 0 6
1471 1494
1512 1494
1512 1383
1128 1383
1128 1452
1182 1452
10 5 9 0 0 0 0 361 361 0 0 6
1477 1467
1484 1467
1484 1409
1373 1409
1373 1485
1407 1485
9 6 127 0 0 12416 0 361 361 0 0 6
1471 1458
1493 1458
1493 1400
1364 1400
1364 1494
1407 1494
12 1 128 0 0 12416 0 362 361 0 0 4
1252 1506
1327 1506
1327 1449
1407 1449
11 2 45 0 0 0 0 362 361 0 0 4
1246 1497
1335 1497
1335 1458
1407 1458
10 6 129 0 0 12416 0 362 362 0 0 6
1252 1470
1271 1470
1271 1401
1146 1401
1146 1497
1182 1497
9 5 26 0 0 0 0 362 362 0 0 6
1246 1461
1263 1461
1263 1410
1155 1410
1155 1488
1182 1488
3 0 124 0 0 0 0 362 0 0 531 5
1176 1470
1175 1470
1175 1432
1398 1432
1398 1468
7 3 124 0 0 0 0 362 362 0 0 4
1176 1506
1175 1506
1175 1470
1176 1470
8 8 125 0 0 12416 0 362 361 0 0 6
1176 1515
1168 1515
1168 1528
1390 1528
1390 1512
1401 1512
8 4 125 0 0 0 0 361 361 0 0 4
1401 1512
1390 1512
1390 1476
1401 1476
4 8 125 0 0 0 0 362 362 0 0 4
1176 1479
1168 1479
1168 1515
1176 1515
11 1 45 0 0 20608 0 362 356 0 0 6
1246 1497
1291 1497
1291 1608
809 1608
809 1712
2273 1712
11 1 10 0 0 20480 0 361 358 0 0 6
1471 1494
1512 1494
1512 1588
786 1588
786 1654
2272 1654
10 1 9 0 0 0 0 361 359 0 0 6
1477 1467
1484 1467
1484 1579
776 1579
776 1627
2272 1627
1 0 124 0 0 0 0 360 0 0 410 2
1025 1452
1025 1470
7 3 124 0 0 0 0 361 361 0 0 4
1401 1503
1398 1503
1398 1467
1401 1467
1 0 124 0 0 0 3 363 0 0 533 2
221 50
221 67
0 3 124 0 0 0 3 0 364 262 0 4
279 67
221 67
221 64
182 64
14 0 47 0 0 8320 0 381 0 0 143 5
503 1227
510 1227
510 1759
763 1759
763 1860
13 0 50 0 0 8320 0 381 0 0 142 5
503 1218
519 1218
519 1775
754 1775
754 1869
12 0 49 0 0 8320 0 381 0 0 0 3
503 1209
528 1209
528 1666
11 0 48 0 0 8320 0 381 0 0 0 3
503 1200
537 1200
537 1528
8 0 81 0 0 0 0 366 0 0 0 4
361 263
335 263
335 161
456 161
7 0 82 0 0 0 0 366 0 0 0 4
361 254
327 254
327 154
457 154
6 0 83 0 0 0 0 366 0 0 0 4
361 245
318 245
318 146
459 146
5 0 61 0 0 0 0 366 0 0 0 4
361 236
309 236
309 138
461 138
1 0 9 0 0 0 0 365 0 0 0 5
526 214
515 214
515 108
50 108
50 109
4 1 130 0 0 4224 0 366 23 0 0 4
361 227
261 227
261 262
260 262
1 0 10 0 0 4224 0 346 0 0 0 2
57 2705
57 319
1 0 11 0 0 4224 0 347 0 0 0 2
86 2647
86 732
1 0 4 0 0 4224 0 335 0 0 0 3
2761 3106
2761 108
1853 108
1 0 8 0 0 4224 0 344 0 0 0 3
2464 2322
2464 814
2098 814
1 0 6 0 0 0 0 343 0 0 0 3
2522 2482
2522 476
2056 476
1 0 7 0 0 0 0 342 0 0 0 4
2576 2761
2551 2761
2551 467
2080 467
1 0 6 0 0 0 0 340 0 0 164 5
2611 2716
2611 449
2017 449
2017 433
1856 433
14 0 6 0 0 0 0 371 0 0 0 5
1217 458
1204 458
1204 381
1716 381
1716 382
13 0 7 0 0 0 0 371 0 0 0 5
1217 449
1213 449
1213 401
1716 401
1716 402
0 0 124 0 0 0 3 0 0 626 253 2
278 1077
278 321
0 0 124 0 0 0 3 0 0 556 0 2
1146 67
725 67
0 4 124 0 0 0 3 0 390 556 0 5
1417 564
1417 797
1176 797
1176 897
1223 897
4 4 124 0 0 0 3 368 372 0 0 8
1221 188
1146 188
1146 67
1417 67
1417 564
1175 564
1175 713
1240 713
12 0 81 0 0 0 0 370 0 0 685 2
1073 548
1013 548
11 0 82 0 0 0 0 370 0 0 684 2
1073 530
984 530
10 0 83 0 0 0 0 370 0 0 686 2
1073 512
954 512
9 0 61 0 0 0 0 370 0 0 687 2
1073 494
924 494
8 0 81 0 0 0 0 390 0 0 685 2
1223 933
1013 933
7 0 82 0 0 0 0 390 0 0 684 2
1223 924
984 924
6 0 83 0 0 0 0 390 0 0 686 2
1223 915
954 915
5 0 61 0 0 0 0 390 0 0 687 2
1223 906
924 906
14 1 131 0 0 4224 0 390 386 0 0 4
1287 933
1444 933
1444 896
1443 896
13 1 132 0 0 4224 0 390 385 0 0 3
1287 924
1420 924
1420 896
12 1 133 0 0 4224 0 390 387 0 0 3
1287 915
1397 915
1397 896
11 1 134 0 0 4224 0 390 388 0 0 3
1287 906
1374 906
1374 896
9 1 2 0 0 0 0 390 389 0 0 2
1293 870
1293 846
3 2 84 0 0 0 0 390 390 0 0 2
1217 888
1217 879
10 9 2 0 0 0 0 390 390 0 0 2
1293 879
1293 870
1 9 2 0 0 0 0 390 390 0 0 5
1223 870
1213 870
1213 850
1293 850
1293 870
8 0 81 0 0 0 0 368 0 0 685 2
1221 224
1013 224
7 0 82 0 0 0 0 368 0 0 684 2
1221 215
984 215
6 0 83 0 0 0 0 368 0 0 686 2
1221 206
954 206
5 0 61 0 0 0 0 368 0 0 687 2
1221 197
924 197
10 1 2 0 0 0 0 368 374 0 0 4
1291 170
1301 170
1301 170
1298 170
3 2 4 0 0 0 0 368 368 0 0 2
1215 179
1215 170
10 9 2 0 0 0 0 368 368 0 0 2
1291 170
1291 161
1 9 2 0 0 0 0 368 368 0 0 5
1221 161
1220 161
1220 141
1291 141
1291 161
12 0 81 0 0 0 0 369 0 0 685 2
1071 345
1013 345
11 0 82 0 0 0 0 369 0 0 684 2
1071 327
984 327
10 0 83 0 0 0 0 369 0 0 686 2
1071 309
954 309
9 0 61 0 0 0 0 369 0 0 687 2
1071 291
924 291
8 0 81 0 0 0 0 384 0 0 685 4
643 1113
618 1113
618 1161
1013 1161
7 0 82 0 0 0 0 384 0 0 684 4
643 1104
609 1104
609 1152
984 1152
6 0 83 0 0 0 0 384 0 0 686 4
643 1095
600 1095
600 1143
954 1143
5 0 61 0 0 0 0 384 0 0 687 4
643 1086
591 1086
591 1134
924 1134
8 0 85 0 0 12288 0 381 0 0 688 4
439 1227
418 1227
418 1277
867 1277
7 0 86 0 0 12288 0 381 0 0 689 4
439 1218
407 1218
407 1267
836 1267
6 0 87 0 0 12288 0 381 0 0 690 4
439 1209
397 1209
397 1258
804 1258
5 0 88 0 0 12288 0 381 0 0 691 4
439 1200
387 1200
387 1248
772 1248
18 0 81 0 0 0 0 378 0 0 252 2
690 711
794 711
17 0 82 0 0 0 0 378 0 0 251 2
690 702
792 702
16 0 83 0 0 0 0 378 0 0 250 2
690 693
793 693
15 0 61 0 0 0 0 378 0 0 0 2
690 684
783 684
14 0 85 0 0 0 0 378 0 0 238 2
690 675
867 675
13 0 86 0 0 0 0 378 0 0 239 2
690 666
836 666
12 0 87 0 0 0 0 378 0 0 240 2
690 657
804 657
11 0 88 0 0 0 0 378 0 0 241 2
690 648
772 648
8 0 81 0 0 0 0 367 0 0 685 4
632 324
650 324
650 350
1013 350
7 0 82 0 0 0 0 367 0 0 684 5
623 324
623 319
657 319
657 332
984 332
6 0 83 0 0 0 0 367 0 0 686 3
614 324
614 312
954 312
5 0 61 0 0 0 0 367 0 0 687 3
605 324
605 297
924 297
12 0 81 0 0 0 0 365 0 0 685 2
590 277
1013 277
11 0 82 0 0 0 0 365 0 0 684 2
590 259
984 259
10 0 83 0 0 0 0 365 0 0 686 2
590 241
954 241
9 0 61 0 0 0 0 365 0 0 687 2
590 223
924 223
2 14 98 0 0 4224 0 376 367 0 0 4
617 490
617 432
632 432
632 388
4 13 99 0 0 4224 0 376 367 0 0 4
599 490
599 423
623 423
623 388
6 12 100 0 0 4224 0 376 367 0 0 4
581 490
581 414
614 414
614 388
8 11 101 0 0 4224 0 376 367 0 0 4
563 490
563 405
605 405
605 388
4 0 124 0 0 0 3 367 0 0 0 4
596 324
596 297
278 297
278 261
2 3 12 0 0 0 0 367 367 0 0 2
578 318
587 318
1 1 2 0 0 0 0 367 373 0 0 3
569 324
569 323
541 323
1 9 2 0 0 0 0 367 367 0 0 5
569 324
569 323
546 323
546 394
569 394
10 9 2 0 0 0 0 367 367 0 0 2
578 394
569 394
14 0 81 0 0 0 0 384 0 0 685 2
707 1113
1013 1113
13 0 82 0 0 0 0 384 0 0 684 2
707 1104
984 1104
12 0 83 0 0 0 0 384 0 0 686 2
707 1095
954 1095
11 0 61 0 0 0 0 384 0 0 687 2
707 1086
924 1086
1 1 2 0 0 0 0 384 383 0 0 3
643 1050
627 1050
627 1044
3 2 15 0 0 0 0 384 381 0 0 5
637 1068
637 1059
422 1059
422 1173
433 1173
3 2 15 0 0 0 0 384 384 0 0 2
637 1068
637 1059
10 9 14 0 0 0 0 384 384 0 0 4
713 1059
714 1059
714 1050
713 1050
4 4 124 0 0 0 3 384 381 0 0 4
643 1077
278 1077
278 1191
439 1191
9 1 2 0 0 0 0 381 382 0 0 4
509 1164
524 1164
524 1164
519 1164
3 2 15 0 0 0 0 381 381 0 0 4
433 1182
422 1182
422 1173
433 1173
10 9 2 0 0 0 0 381 381 0 0 4
509 1173
510 1173
510 1164
509 1164
1 9 2 0 0 0 0 381 381 0 0 6
439 1164
438 1164
438 1144
510 1144
510 1164
509 1164
1 1 135 0 0 8320 0 36 379 0 0 4
610 919
610 908
743 908
743 816
10 1 2 0 0 0 0 379 380 0 0 5
662 822
662 826
641 826
641 795
633 795
3 1 112 0 0 8320 0 379 33 0 0 4
725 816
725 859
540 859
540 898
5 1 113 0 0 8320 0 379 32 0 0 4
707 816
707 850
512 850
512 897
7 1 114 0 0 8320 0 379 34 0 0 4
689 816
689 840
484 840
484 897
9 1 115 0 0 8320 0 379 35 0 0 4
671 816
671 831
452 831
452 897
2 0 81 0 0 0 0 379 0 0 685 3
734 816
734 859
1013 859
4 0 82 0 0 0 0 379 0 0 684 3
716 816
716 849
984 849
6 0 83 0 0 0 0 379 0 0 686 3
698 816
698 840
954 840
8 0 61 0 0 0 0 379 0 0 687 3
680 816
680 831
924 831
13 0 111 0 0 4224 0 379 0 0 0 4
689 752
689 736
702 736
702 722
14 0 110 0 0 4224 0 379 0 0 0 4
671 752
671 725
697 725
697 719
10 11 106 0 0 8320 0 378 376 0 0 3
626 711
608 711
608 554
9 12 107 0 0 8320 0 378 376 0 0 3
626 702
590 702
590 554
8 13 108 0 0 8320 0 378 376 0 0 3
626 693
572 693
572 554
7 14 109 0 0 8320 0 378 376 0 0 3
626 684
554 684
554 554
19 1 13 0 0 0 0 378 322 0 0 6
696 630
700 630
700 600
511 600
511 673
174 673
1 1 136 0 0 8320 0 376 31 0 0 3
626 490
626 459
669 459
1 3 102 0 0 8320 0 28 376 0 0 4
462 510
462 471
608 471
608 490
1 5 103 0 0 8320 0 27 376 0 0 4
434 510
434 461
590 461
590 490
1 7 104 0 0 8320 0 29 376 0 0 4
405 510
405 451
572 451
572 490
1 9 105 0 0 8320 0 30 376 0 0 4
374 510
374 442
554 442
554 490
1 10 2 0 0 0 0 377 376 0 0 3
528 504
528 484
545 484
9 1 2 0 0 0 0 372 375 0 0 5
1310 686
1291 686
1291 617
1284 617
1284 613
3 2 19 0 0 0 0 372 372 0 0 7
1234 704
1224 704
1224 650
1216 650
1216 650
1234 650
1234 695
10 9 2 0 0 0 0 372 372 0 0 4
1310 695
1310 641
1310 641
1310 686
1 9 2 0 0 0 0 372 372 0 0 5
1240 686
1212 686
1212 617
1310 617
1310 686
0 8 116 0 0 4096 0 0 371 669 0 3
1349 345
1349 512
1287 512
0 7 117 0 0 4096 0 0 371 670 0 3
1335 327
1335 503
1287 503
0 6 118 0 0 4096 0 0 371 671 0 3
1321 309
1321 494
1287 494
0 5 119 0 0 4224 0 0 371 672 0 3
1308 291
1308 485
1287 485
8 22 120 0 0 4224 0 370 371 0 0 2
1137 548
1211 548
6 21 121 0 0 4224 0 370 371 0 0 4
1137 530
1184 530
1184 539
1211 539
20 4 122 0 0 12416 0 371 370 0 0 4
1211 530
1195 530
1195 512
1137 512
2 19 123 0 0 4224 0 370 371 0 0 4
1137 494
1206 494
1206 521
1211 521
5 7 2 0 0 0 0 370 370 0 0 4
1137 521
1166 521
1166 539
1137 539
3 5 2 0 0 0 0 370 370 0 0 4
1137 503
1166 503
1166 521
1137 521
1 3 2 0 0 0 0 370 370 0 0 4
1137 485
1166 485
1166 503
1137 503
8 14 116 0 0 4224 0 369 368 0 0 4
1135 345
1349 345
1349 224
1285 224
6 13 117 0 0 4224 0 369 368 0 0 4
1135 327
1335 327
1335 215
1285 215
4 12 118 0 0 4224 0 369 368 0 0 4
1135 309
1321 309
1321 206
1285 206
2 11 119 0 0 0 0 369 368 0 0 4
1135 291
1308 291
1308 197
1285 197
1 0 5 0 0 0 0 369 0 0 0 4
1135 282
1144 282
1144 270
1725 270
5 7 5 0 0 0 0 369 369 0 0 4
1135 318
1144 318
1144 336
1135 336
3 5 5 0 0 0 0 369 369 0 0 4
1135 300
1144 300
1144 318
1135 318
1 3 5 0 0 0 0 369 369 0 0 4
1135 282
1144 282
1144 300
1135 300
11 2 97 0 0 12416 0 366 365 0 0 4
425 236
458 236
458 223
526 223
14 8 94 0 0 12416 0 366 365 0 0 4
425 263
457 263
457 277
526 277
13 6 95 0 0 12416 0 366 365 0 0 4
425 254
468 254
468 259
526 259
12 4 96 0 0 12416 0 366 365 0 0 4
425 245
468 245
468 241
526 241
7 5 9 0 0 0 0 365 365 0 0 4
526 268
515 268
515 250
526 250
5 3 9 0 0 0 0 365 365 0 0 4
526 250
515 250
515 232
526 232
3 1 9 0 0 0 0 365 365 0 0 4
526 232
515 232
515 214
526 214
0 0 82 0 0 4224 0 0 0 0 0 2
984 1369
984 128
0 1 81 0 0 4224 0 0 0 0 0 2
1013 1369
1013 126
0 0 83 0 0 4224 0 0 0 0 0 2
954 1369
954 129
0 0 61 0 0 4224 0 0 0 0 0 2
924 1369
924 130
0 0 85 0 0 4224 0 0 0 0 0 2
867 1369
867 782
0 0 86 0 0 4224 0 0 0 0 0 2
836 1369
836 783
0 0 87 0 0 4224 0 0 0 0 0 2
804 1369
804 784
0 0 88 0 0 4224 0 0 0 0 0 2
772 1369
772 784
256
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1450 493 1520 508
1464 504 1505 515
6 lb Bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2826 766 2896 781
2840 777 2881 788
6 lb Bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
526 18 615 39
534 25 606 40
9 CLK PULSE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
2271 1737 2380 1761
2281 1745 2369 1761
11 LDAM (0000)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1515 545 1584 569
1525 553 1573 569
6 Lc BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1572 781 1617 805
1582 789 1606 805
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 2460 45 2484
21 2465 37 2481
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 2402 75 2426
51 2407 67 2423
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
61 2348 124 2372
68 2354 116 2370
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
89 2286 152 2310
96 2292 144 2308
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
143 2189 206 2213
150 2195 198 2211
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
199 2050 262 2074
206 2056 254 2072
6 Li BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
169 2002 232 2026
176 2007 224 2023
6 Ei BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
143 1953 206 1977
150 1959 198 1975
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
88 1838 151 1862
95 1844 143 1860
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
59 1783 122 1807
66 1789 114 1805
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
43 1739 74 1763
50 1744 66 1760
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 1701 45 1725
21 1706 37 1722
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 1137 45 1161
21 1142 37 1158
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
43 1178 74 1202
50 1183 66 1199
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
59 1218 122 1242
66 1224 114 1240
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
88 1252 151 1276
95 1258 143 1274
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 722 45 746
21 727 37 743
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 746 75 770
51 751 67 767
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 414 45 438
21 419 37 435
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 447 75 471
51 452 67 468
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
58 782 121 806
65 788 113 804
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
59 486 122 510
66 492 114 508
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
86 829 149 853
93 835 141 851
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
88 525 151 549
95 531 143 547
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
143 1334 206 1358
150 1340 198 1356
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
143 909 206 933
150 915 198 931
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
169 1382 232 1406
176 1387 224 1403
6 Ei BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
197 1437 260 1461
204 1443 252 1459
6 Li BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2434 2153 2497 2177
2441 2158 2489 2174
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2435 1877 2498 1901
2442 1882 2490 1898
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2434 1548 2497 1572
2441 1553 2489 1569
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2433 1215 2496 1239
2440 1220 2488 1236
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2433 947 2496 971
2440 952 2488 968
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 2425 2599 2446
2574 2432 2590 2447
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2596 2462 2627 2486
2603 2468 2619 2484
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2624 2511 2663 2535
2631 2517 2655 2533
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 2597 2683 2621
2667 2603 2675 2619
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2716 2723 2747 2747
2723 2729 2739 2745
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2736 2795 2799 2819
2743 2800 2791 2816
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2737 2374 2800 2398
2744 2379 2792 2395
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2738 2081 2801 2105
2745 2086 2793 2102
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 2351 2748 2375
2724 2357 2740 2373
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 2061 2748 2085
2724 2067 2740 2083
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2689 2331 2720 2355
2696 2336 2712 2352
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2689 2041 2720 2065
2696 2046 2712 2062
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 2312 2683 2336
2667 2318 2675 2334
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 2022 2683 2046
2667 2028 2675 2044
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 2292 2664 2316
2632 2298 2656 2314
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 2004 2664 2028
2632 2010 2656 2026
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2596 2276 2627 2300
2603 2282 2619 2298
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2596 1988 2627 2012
2603 1994 2619 2010
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 2258 2599 2279
2574 2265 2590 2280
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 1971 2599 1992
2574 1978 2590 1993
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2738 1743 2801 1767
2745 1748 2793 1764
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 1723 2748 1747
2724 1729 2740 1745
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 1693 2683 1717
2667 1699 2675 1715
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2738 1412 2801 1436
2745 1417 2793 1433
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2737 1139 2800 1163
2744 1144 2792 1160
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 1392 2748 1416
2724 1398 2740 1414
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 1124 2748 1148
2724 1130 2740 1146
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2736 913 2799 937
2743 918 2791 934
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 893 2748 917
2724 899 2740 915
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 1362 2683 1386
2667 1368 2675 1384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 1098 2683 1122
2667 1104 2675 1120
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 1677 2664 1701
2632 1683 2656 1699
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2596 1663 2627 1687
2603 1669 2619 1685
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2565 1648 2598 1669
2573 1655 2589 1670
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 1348 2664 1372
2632 1354 2656 1370
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2596 1336 2627 1360
2603 1342 2619 1358
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 1319 2599 1340
2574 1326 2590 1341
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 1086 2664 1110
2632 1092 2656 1108
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 859 2683 883
2667 865 2675 881
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 837 2664 861
2632 843 2656 859
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2595 1069 2626 1093
2602 1075 2618 1091
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 1052 2597 1076
2573 1058 2589 1074
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2595 809 2626 833
2602 815 2618 831
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2736 510 2799 534
2743 515 2791 531
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2737 290 2800 314
2744 295 2792 311
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2717 486 2748 510
2724 492 2740 508
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2567 789 2598 813
2574 795 2590 811
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2537 2238 2568 2262
2544 2244 2560 2260
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2536 1952 2567 1976
2543 1958 2559 1974
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2536 1632 2567 1656
2543 1638 2559 1654
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2536 1303 2567 1327
2543 1309 2559 1325
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2536 1036 2567 1060
2543 1042 2559 1058
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2537 767 2568 791
2544 773 2560 789
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2507 2219 2538 2243
2514 2225 2530 2241
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1932 2537 1956
2513 1938 2529 1954
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1612 2537 1636
2513 1618 2529 1634
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1284 2537 1308
2513 1290 2529 1306
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 1017 2537 1041
2513 1023 2529 1039
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2507 743 2538 767
2514 749 2530 765
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2705 89 2768 113
2712 94 2760 110
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2371 88 2434 112
2378 93 2426 109
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1932 89 1995 113
1939 94 1987 110
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2708 249 2739 273
2715 255 2731 271
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2368 250 2399 274
2375 256 2391 272
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1945 249 1976 273
1952 255 1968 271
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1208 394 1247 418
1215 400 1239 416
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1190 377 1213 401
1197 383 1205 399
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2660 436 2683 460
2667 442 2675 458
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2625 414 2664 438
2632 420 2656 436
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2293 382 2332 406
2300 388 2324 404
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2332 362 2355 386
2339 368 2347 384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1953 362 1976 386
1960 368 1968 384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1911 382 1950 406
1918 388 1942 404
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2078 436 2109 460
2085 442 2101 458
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2114 444 2145 468
2121 450 2137 466
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2146 453 2177 477
2153 459 2169 475
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2178 462 2209 486
2185 468 2201 484
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2597 513 2628 537
2604 519 2620 535
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2566 498 2597 522
2573 504 2589 520
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1736 435 1767 459
1743 441 1759 457
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1763 444 1794 468
1770 450 1786 466
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1816 462 1847 486
1823 468 1839 484
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1787 453 1818 477
1794 459 1810 475
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2537 482 2568 506
2544 488 2560 504
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2506 473 2537 497
2513 479 2529 495
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2378 787 2441 811
2385 792 2433 808
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2303 1616 2334 1640
2310 1621 2326 1637
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2305 1646 2336 1670
2312 1651 2328 1667
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2306 1672 2337 1696
2313 1678 2329 1694
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2306 1699 2337 1723
2313 1705 2329 1721
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
818 1690 849 1714
825 1696 841 1712
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
818 1661 849 1685
825 1667 841 1683
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
817 1634 848 1658
824 1639 840 1655
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
818 1608 849 1632
825 1613 841 1629
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1346 842 1473 866
1353 847 1465 863
14 BINARY DISPLAY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1214 817 1285 841
1221 822 1277 838
7 O/P REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
552 1191 763 1215
557 1195 757 1211
25 8 bit From RAM  <<<---<<<
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
583 1161 754 1185
588 1165 748 1181
20 LSB 4 BIT -> address
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
583 1226 746 1250
588 1230 740 1246
19 MSB 4 BIT -> opcode
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
938 89 993 113
945 94 985 110
5 VALUE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
785 89 856 113
792 94 848 110
7 ADDRESS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
524 162 623 186
529 166 617 182
11 BUFFER-> PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
380 161 407 185
385 165 401 181
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
642 343 677 367
647 347 671 363
3 MAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1235 114 1270 138
1240 118 1264 134
3 ACC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1050 245 1157 269
1055 249 1151 265
12 BUFFER-> ACC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1232 410 1275 431
1241 416 1265 431
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1042 445 1149 469
1047 449 1143 465
12 BUFFER-> ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
938 108 969 132
945 113 961 129
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
969 107 1000 131
976 113 992 129
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
999 107 1030 131
1006 113 1022 129
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
757 108 788 132
764 114 780 130
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 109 819 133
795 114 811 130
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
820 109 851 133
827 114 843 130
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
852 108 883 132
859 113 875 129
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
640 510 679 534
647 515 671 531
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
357 549 388 573
364 554 380 570
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
390 548 421 572
397 554 413 570
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
419 549 450 573
426 554 442 570
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
449 548 480 572
456 554 472 570
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
365 571 476 615
372 577 468 609
23 Address From 
    USER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
639 563 678 587
646 569 670 585
3 RAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
442 947 537 991
449 952 529 984
21 Value From 
    USER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
436 930 467 954
443 935 459 951
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
468 929 499 953
475 935 491 951
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
498 931 529 955
505 936 521 952
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
527 930 558 954
534 936 550 952
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
596 939 627 963
603 945 619 961
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
689 446 720 470
696 451 712 467
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
442 1089 505 1153
449 1095 497 1143
18   IR
 MSB
OPCODE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
639 961 710 1025
646 966 702 1014
19   IR
 LSB
ADDRESS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
556 764 595 788
563 769 587 785
3 MUX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1367 44 1406 68
1374 49 1398 65
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1378 539 1417 563
1385 544 1409 560
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1376 769 1415 793
1383 774 1407 790
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
275 64 314 88
282 69 306 85
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
274 274 313 298
281 279 305 295
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
878 43 917 67
885 48 909 64
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
272 1053 311 1077
279 1058 303 1074
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
277 1168 316 1192
284 1173 308 1189
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
200 280 263 304
207 286 255 302
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
208 617 271 641
215 623 263 639
6 WE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
208 647 271 671
215 653 263 669
6 CE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
217 996 280 1020
224 1001 272 1017
6 Ei BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
213 1143 276 1167
220 1149 268 1165
6 Li BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1509 87 1572 111
1516 92 1564 108
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1490 362 1513 386
1497 368 1505 384
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1452 382 1491 406
1459 388 1483 404
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 433 1478 457
1454 439 1470 455
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 442 1478 466
1454 448 1470 464
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 452 1478 476
1454 458 1470 474
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1447 462 1478 486
1454 468 1470 484
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1454 788 1517 812
1461 793 1509 809
6 Lo BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
273 875 312 899
280 880 304 896
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1513 249 1544 273
1520 255 1536 271
2 Ea
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
1510 322 1559 370
1517 327 1551 359
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
216 190 247 214
223 195 239 211
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
226 85 257 109
233 90 249 106
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
482 84 513 108
489 89 505 105
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1140 366 1171 390
1147 371 1163 387
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1164 247 1195 271
1171 253 1187 269
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
116 29 205 50
124 36 196 51
9 CLK PULSE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1508 1531 1539 1555
1515 1536 1531 1552
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1239 1541 1270 1565
1246 1547 1262 1563
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1288 1541 1319 1565
1295 1547 1311 1563
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1270 1337 1381 1361
1277 1342 1373 1358
12 RING COUNTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1535 1426 1574 1470
1542 1431 1566 1463
7 F/F
 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1537 1475 1576 1519
1544 1481 1568 1513
7 F/F
 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1078 1429 1117 1473
1085 1435 1109 1467
7 F/F
 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1108 1475 1147 1519
1115 1480 1139 1512
7 F/F
 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
472 1405 575 1429
479 1411 567 1427
11 I4 I5 I6 I7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1162 105 1225 129
1169 110 1217 126
6 La BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
434 296 497 320
441 302 489 318
6 Lm BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
701 592 764 616
708 598 756 614
6 WE BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
274 412 313 436
281 417 305 433
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
795 1470 882 1494
802 1476 874 1492
9 CLK PULSE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
278 1444 317 1468
285 1449 309 1465
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
670 1446 709 1470
677 1451 701 1467
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
946 1447 985 1471
953 1452 977 1468
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
201 210 264 234
208 216 256 232
6 Lp BAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
3082 598 3119 622
3092 606 3108 622
2 ZF
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
3078 1076 3115 1100
3088 1084 3104 1100
2 ZF
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
3086 1468 3123 1492
3096 1476 3112 1492
2 ZF
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1489 1284 1616 1306
1496 1292 1608 1308
14 CONTROL MATRIX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
876 1509 969 1533
886 1517 958 1533
9 For Check
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
416 282 455 306
423 287 447 303
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
97 236 240 280
104 242 232 274
29 0 -> CLR (Reset)
1 -> Active
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
46 107 136 130
59 117 122 132
9 EP SNIPED
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
911 105 944 129
919 113 935 129
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1807 563 1868 587
1817 571 1857 587
5 C REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1215 586 1276 610
1225 594 1265 610
5 B REG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1837 986 1870 1010
1845 994 1861 1010
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1849 849 1882 873
1857 857 1873 873
2 C3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1118 770 1151 794
1126 778 1142 794
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1116 654 1149 678
1124 662 1140 678
2 B3
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
306 732 417 758
316 740 406 758
9 SIGN FLAG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
1036 1535 1185 1579
1046 1543 1174 1575
29 1 -> CLR (Reset)
0 -> Active
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
359 1896 476 1920
369 1904 465 1920
12 control unit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1060 2133 1097 2157
1070 2141 1086 2157
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1150 2298 1219 2322
1160 2306 1208 2322
6 lm bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1229 2270 1272 2285
1243 2281 1257 2292
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1319 2259 1389 2274
1333 2270 1374 2281
6 Li bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1649 2367 1719 2382
1663 2379 1704 2390
6 sub t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1761 2369 1828 2384
1776 2380 1812 2391
5 xr t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1669 2610 1739 2625
1683 2621 1724 2632
6 la bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1800 2631 1870 2646
1814 2643 1855 2654
6 Ei bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1940 2630 2010 2645
1954 2641 1995 2652
6 lb bar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2066 2636 2109 2651
2080 2647 2094 2658
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2176 2601 2219 2616
2190 2613 2204 2624
2 Lo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1882 2429 1949 2444
1897 2440 1933 2451
5 Jz t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2207 2723 2301 2738
2222 2734 2285 2745
9 s1 s2 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
2316 2527 2394 2542
2330 2539 2379 2550
7 Se S3 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2414 2599 2459 2614
2429 2610 2443 2621
2 Zf
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2480 2636 2523 2651
2494 2647 2508 2658
2 Lp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
1464 2349 1492 2416
1474 2359 1481 2414
18 C
e 
b
a
r
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1153 2118 1222 2142
1163 2126 1211 2142
6 lda t3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1086 1802 1111 1846
1094 1810 1102 1842
5 T
1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
